`timescale 1 ns/100 ps
// Version: 2022.1 2022.1.0.10


module PF_DRI_C0_PF_DRI_C0_0_PF_DRI(
       PCLK,
       PSEL,
       PENABLE,
       PWRITE,
       PADDR,
       PSTRB,
       PWDATA,
       PRESETN,
       PRDATA,
       PREADY,
       PSLVERR,
       PINTERRUPT,
       PTIMEOUT,
       BUSERROR,
       Q0_LANE0_DRI_CTRL,
       Q0_LANE0_DRI_RDATA,
       Q0_LANE0_DRI_INTERRUPT,
       Q0_LANE1_DRI_CTRL,
       Q0_LANE1_DRI_RDATA,
       Q0_LANE1_DRI_INTERRUPT,
       Q0_LANE2_DRI_CTRL,
       Q0_LANE2_DRI_RDATA,
       Q0_LANE2_DRI_INTERRUPT,
       Q0_LANE3_DRI_CTRL,
       Q0_LANE3_DRI_RDATA,
       Q0_LANE3_DRI_INTERRUPT,
       Q1_LANE0_DRI_CTRL,
       Q1_LANE0_DRI_RDATA,
       Q1_LANE0_DRI_INTERRUPT,
       Q1_LANE1_DRI_CTRL,
       Q1_LANE1_DRI_RDATA,
       Q1_LANE1_DRI_INTERRUPT,
       Q1_LANE2_DRI_CTRL,
       Q1_LANE2_DRI_RDATA,
       Q1_LANE2_DRI_INTERRUPT,
       Q1_LANE3_DRI_CTRL,
       Q1_LANE3_DRI_RDATA,
       Q1_LANE3_DRI_INTERRUPT,
       Q2_LANE0_DRI_CTRL,
       Q2_LANE0_DRI_RDATA,
       Q2_LANE0_DRI_INTERRUPT,
       Q2_LANE1_DRI_CTRL,
       Q2_LANE1_DRI_RDATA,
       Q2_LANE1_DRI_INTERRUPT,
       Q2_LANE2_DRI_CTRL,
       Q2_LANE2_DRI_RDATA,
       Q2_LANE2_DRI_INTERRUPT,
       Q2_LANE3_DRI_CTRL,
       Q2_LANE3_DRI_RDATA,
       Q2_LANE3_DRI_INTERRUPT,
       Q3_LANE0_DRI_CTRL,
       Q3_LANE0_DRI_RDATA,
       Q3_LANE0_DRI_INTERRUPT,
       Q3_LANE1_DRI_CTRL,
       Q3_LANE1_DRI_RDATA,
       Q3_LANE1_DRI_INTERRUPT,
       Q3_LANE2_DRI_CTRL,
       Q3_LANE2_DRI_RDATA,
       Q3_LANE2_DRI_INTERRUPT,
       Q3_LANE3_DRI_CTRL,
       Q3_LANE3_DRI_RDATA,
       Q3_LANE3_DRI_INTERRUPT,
       Q4_LANE0_DRI_CTRL,
       Q4_LANE0_DRI_RDATA,
       Q4_LANE0_DRI_INTERRUPT,
       Q4_LANE1_DRI_CTRL,
       Q4_LANE1_DRI_RDATA,
       Q4_LANE1_DRI_INTERRUPT,
       Q4_LANE2_DRI_CTRL,
       Q4_LANE2_DRI_RDATA,
       Q4_LANE2_DRI_INTERRUPT,
       Q4_LANE3_DRI_CTRL,
       Q4_LANE3_DRI_RDATA,
       Q4_LANE3_DRI_INTERRUPT,
       Q5_LANE0_DRI_CTRL,
       Q5_LANE0_DRI_RDATA,
       Q5_LANE0_DRI_INTERRUPT,
       Q5_LANE1_DRI_CTRL,
       Q5_LANE1_DRI_RDATA,
       Q5_LANE1_DRI_INTERRUPT,
       Q5_LANE2_DRI_CTRL,
       Q5_LANE2_DRI_RDATA,
       Q5_LANE2_DRI_INTERRUPT,
       Q5_LANE3_DRI_CTRL,
       Q5_LANE3_DRI_RDATA,
       Q5_LANE3_DRI_INTERRUPT,
       Q4_TXPLL_SSC_DRI_CTRL,
       Q4_TXPLL_SSC_DRI_RDATA,
       Q4_TXPLL_SSC_DRI_INTERRUPT,
       Q2_TXPLL_SSC_DRI_CTRL,
       Q2_TXPLL_SSC_DRI_RDATA,
       Q2_TXPLL_SSC_DRI_INTERRUPT,
       Q0_TXPLL_SSC_DRI_CTRL,
       Q0_TXPLL_SSC_DRI_RDATA,
       Q0_TXPLL_SSC_DRI_INTERRUPT,
       Q1_TXPLL_SSC_DRI_CTRL,
       Q1_TXPLL_SSC_DRI_RDATA,
       Q1_TXPLL_SSC_DRI_INTERRUPT,
       Q3_TXPLL_SSC_DRI_CTRL,
       Q3_TXPLL_SSC_DRI_RDATA,
       Q3_TXPLL_SSC_DRI_INTERRUPT,
       Q5_TXPLL_SSC_DRI_CTRL,
       Q5_TXPLL_SSC_DRI_RDATA,
       Q5_TXPLL_SSC_DRI_INTERRUPT,
       Q4_TXPLL_DRI_CTRL,
       Q4_TXPLL_DRI_RDATA,
       Q4_TXPLL_DRI_INTERRUPT,
       Q2_TXPLL0_DRI_CTRL,
       Q2_TXPLL0_DRI_RDATA,
       Q2_TXPLL0_DRI_INTERRUPT,
       Q2_TXPLL1_DRI_CTRL,
       Q2_TXPLL1_DRI_RDATA,
       Q2_TXPLL1_DRI_INTERRUPT,
       Q0_TXPLL0_DRI_CTRL,
       Q0_TXPLL0_DRI_RDATA,
       Q0_TXPLL0_DRI_INTERRUPT,
       Q0_TXPLL1_DRI_CTRL,
       Q0_TXPLL1_DRI_RDATA,
       Q0_TXPLL1_DRI_INTERRUPT,
       Q1_TXPLL0_DRI_CTRL,
       Q1_TXPLL0_DRI_RDATA,
       Q1_TXPLL0_DRI_INTERRUPT,
       Q1_TXPLL1_DRI_CTRL,
       Q1_TXPLL1_DRI_RDATA,
       Q1_TXPLL1_DRI_INTERRUPT,
       Q3_TXPLL_DRI_CTRL,
       Q3_TXPLL_DRI_RDATA,
       Q3_TXPLL_DRI_INTERRUPT,
       Q5_TXPLL_DRI_CTRL,
       Q5_TXPLL_DRI_RDATA,
       Q5_TXPLL_DRI_INTERRUPT,
       PLL0_NW_DRI_CTRL,
       PLL0_NW_DRI_RDATA,
       PLL0_NW_DRI_INTERRUPT,
       PLL1_NW_DRI_CTRL,
       PLL1_NW_DRI_RDATA,
       PLL1_NW_DRI_INTERRUPT,
       PLL0_NE_DRI_CTRL,
       PLL0_NE_DRI_RDATA,
       PLL0_NE_DRI_INTERRUPT,
       PLL1_NE_DRI_CTRL,
       PLL1_NE_DRI_RDATA,
       PLL1_NE_DRI_INTERRUPT,
       PLL0_SE_DRI_CTRL,
       PLL0_SE_DRI_RDATA,
       PLL0_SE_DRI_INTERRUPT,
       PLL1_SE_DRI_CTRL,
       PLL1_SE_DRI_RDATA,
       PLL1_SE_DRI_INTERRUPT,
       PLL0_SW_DRI_CTRL,
       PLL0_SW_DRI_RDATA,
       PLL0_SW_DRI_INTERRUPT,
       PLL1_SW_DRI_CTRL,
       PLL1_SW_DRI_RDATA,
       PLL1_SW_DRI_INTERRUPT,
       DLL0_NW_DRI_CTRL,
       DLL0_NW_DRI_RDATA,
       DLL0_NW_DRI_INTERRUPT,
       DLL1_NW_DRI_CTRL,
       DLL1_NW_DRI_RDATA,
       DLL1_NW_DRI_INTERRUPT,
       DLL0_NE_DRI_CTRL,
       DLL0_NE_DRI_RDATA,
       DLL0_NE_DRI_INTERRUPT,
       DLL1_NE_DRI_CTRL,
       DLL1_NE_DRI_RDATA,
       DLL1_NE_DRI_INTERRUPT,
       DLL0_SE_DRI_CTRL,
       DLL0_SE_DRI_RDATA,
       DLL0_SE_DRI_INTERRUPT,
       DLL1_SE_DRI_CTRL,
       DLL1_SE_DRI_RDATA,
       DLL1_SE_DRI_INTERRUPT,
       DLL0_SW_DRI_CTRL,
       DLL0_SW_DRI_RDATA,
       DLL0_SW_DRI_INTERRUPT,
       DLL1_SW_DRI_CTRL,
       DLL1_SW_DRI_RDATA,
       DLL1_SW_DRI_INTERRUPT,
       CRYPTO_DRI_CTRL,
       CRYPTO_DRI_RDATA,
       CRYPTO_DRI_INTERRUPT,
       DRI_CLK,
       DRI_WDATA,
       DRI_ARST_N
    );
input  PCLK;
input  PSEL;
input  PENABLE;
input  PWRITE;
input  [28:0] PADDR;
input  [3:0] PSTRB;
input  [31:0] PWDATA;
input  PRESETN;
output [31:0] PRDATA;
output PREADY;
output PSLVERR;
output PINTERRUPT;
output PTIMEOUT;
output BUSERROR;
output [10:0] Q0_LANE0_DRI_CTRL;
input  [32:0] Q0_LANE0_DRI_RDATA;
input  Q0_LANE0_DRI_INTERRUPT;
output [10:0] Q0_LANE1_DRI_CTRL;
input  [32:0] Q0_LANE1_DRI_RDATA;
input  Q0_LANE1_DRI_INTERRUPT;
output [10:0] Q0_LANE2_DRI_CTRL;
input  [32:0] Q0_LANE2_DRI_RDATA;
input  Q0_LANE2_DRI_INTERRUPT;
output [10:0] Q0_LANE3_DRI_CTRL;
input  [32:0] Q0_LANE3_DRI_RDATA;
input  Q0_LANE3_DRI_INTERRUPT;
output [10:0] Q1_LANE0_DRI_CTRL;
input  [32:0] Q1_LANE0_DRI_RDATA;
input  Q1_LANE0_DRI_INTERRUPT;
output [10:0] Q1_LANE1_DRI_CTRL;
input  [32:0] Q1_LANE1_DRI_RDATA;
input  Q1_LANE1_DRI_INTERRUPT;
output [10:0] Q1_LANE2_DRI_CTRL;
input  [32:0] Q1_LANE2_DRI_RDATA;
input  Q1_LANE2_DRI_INTERRUPT;
output [10:0] Q1_LANE3_DRI_CTRL;
input  [32:0] Q1_LANE3_DRI_RDATA;
input  Q1_LANE3_DRI_INTERRUPT;
output [10:0] Q2_LANE0_DRI_CTRL;
input  [32:0] Q2_LANE0_DRI_RDATA;
input  Q2_LANE0_DRI_INTERRUPT;
output [10:0] Q2_LANE1_DRI_CTRL;
input  [32:0] Q2_LANE1_DRI_RDATA;
input  Q2_LANE1_DRI_INTERRUPT;
output [10:0] Q2_LANE2_DRI_CTRL;
input  [32:0] Q2_LANE2_DRI_RDATA;
input  Q2_LANE2_DRI_INTERRUPT;
output [10:0] Q2_LANE3_DRI_CTRL;
input  [32:0] Q2_LANE3_DRI_RDATA;
input  Q2_LANE3_DRI_INTERRUPT;
output [10:0] Q3_LANE0_DRI_CTRL;
input  [32:0] Q3_LANE0_DRI_RDATA;
input  Q3_LANE0_DRI_INTERRUPT;
output [10:0] Q3_LANE1_DRI_CTRL;
input  [32:0] Q3_LANE1_DRI_RDATA;
input  Q3_LANE1_DRI_INTERRUPT;
output [10:0] Q3_LANE2_DRI_CTRL;
input  [32:0] Q3_LANE2_DRI_RDATA;
input  Q3_LANE2_DRI_INTERRUPT;
output [10:0] Q3_LANE3_DRI_CTRL;
input  [32:0] Q3_LANE3_DRI_RDATA;
input  Q3_LANE3_DRI_INTERRUPT;
output [10:0] Q4_LANE0_DRI_CTRL;
input  [32:0] Q4_LANE0_DRI_RDATA;
input  Q4_LANE0_DRI_INTERRUPT;
output [10:0] Q4_LANE1_DRI_CTRL;
input  [32:0] Q4_LANE1_DRI_RDATA;
input  Q4_LANE1_DRI_INTERRUPT;
output [10:0] Q4_LANE2_DRI_CTRL;
input  [32:0] Q4_LANE2_DRI_RDATA;
input  Q4_LANE2_DRI_INTERRUPT;
output [10:0] Q4_LANE3_DRI_CTRL;
input  [32:0] Q4_LANE3_DRI_RDATA;
input  Q4_LANE3_DRI_INTERRUPT;
output [10:0] Q5_LANE0_DRI_CTRL;
input  [32:0] Q5_LANE0_DRI_RDATA;
input  Q5_LANE0_DRI_INTERRUPT;
output [10:0] Q5_LANE1_DRI_CTRL;
input  [32:0] Q5_LANE1_DRI_RDATA;
input  Q5_LANE1_DRI_INTERRUPT;
output [10:0] Q5_LANE2_DRI_CTRL;
input  [32:0] Q5_LANE2_DRI_RDATA;
input  Q5_LANE2_DRI_INTERRUPT;
output [10:0] Q5_LANE3_DRI_CTRL;
input  [32:0] Q5_LANE3_DRI_RDATA;
input  Q5_LANE3_DRI_INTERRUPT;
output [10:0] Q4_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q4_TXPLL_SSC_DRI_RDATA;
input  Q4_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q2_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q2_TXPLL_SSC_DRI_RDATA;
input  Q2_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q0_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q0_TXPLL_SSC_DRI_RDATA;
input  Q0_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q1_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q1_TXPLL_SSC_DRI_RDATA;
input  Q1_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q3_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q3_TXPLL_SSC_DRI_RDATA;
input  Q3_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q5_TXPLL_SSC_DRI_CTRL;
input  [32:0] Q5_TXPLL_SSC_DRI_RDATA;
input  Q5_TXPLL_SSC_DRI_INTERRUPT;
output [10:0] Q4_TXPLL_DRI_CTRL;
input  [32:0] Q4_TXPLL_DRI_RDATA;
input  Q4_TXPLL_DRI_INTERRUPT;
output [10:0] Q2_TXPLL0_DRI_CTRL;
input  [32:0] Q2_TXPLL0_DRI_RDATA;
input  Q2_TXPLL0_DRI_INTERRUPT;
output [10:0] Q2_TXPLL1_DRI_CTRL;
input  [32:0] Q2_TXPLL1_DRI_RDATA;
input  Q2_TXPLL1_DRI_INTERRUPT;
output [10:0] Q0_TXPLL0_DRI_CTRL;
input  [32:0] Q0_TXPLL0_DRI_RDATA;
input  Q0_TXPLL0_DRI_INTERRUPT;
output [10:0] Q0_TXPLL1_DRI_CTRL;
input  [32:0] Q0_TXPLL1_DRI_RDATA;
input  Q0_TXPLL1_DRI_INTERRUPT;
output [10:0] Q1_TXPLL0_DRI_CTRL;
input  [32:0] Q1_TXPLL0_DRI_RDATA;
input  Q1_TXPLL0_DRI_INTERRUPT;
output [10:0] Q1_TXPLL1_DRI_CTRL;
input  [32:0] Q1_TXPLL1_DRI_RDATA;
input  Q1_TXPLL1_DRI_INTERRUPT;
output [10:0] Q3_TXPLL_DRI_CTRL;
input  [32:0] Q3_TXPLL_DRI_RDATA;
input  Q3_TXPLL_DRI_INTERRUPT;
output [10:0] Q5_TXPLL_DRI_CTRL;
input  [32:0] Q5_TXPLL_DRI_RDATA;
input  Q5_TXPLL_DRI_INTERRUPT;
output [10:0] PLL0_NW_DRI_CTRL;
input  [32:0] PLL0_NW_DRI_RDATA;
input  PLL0_NW_DRI_INTERRUPT;
output [10:0] PLL1_NW_DRI_CTRL;
input  [32:0] PLL1_NW_DRI_RDATA;
input  PLL1_NW_DRI_INTERRUPT;
output [10:0] PLL0_NE_DRI_CTRL;
input  [32:0] PLL0_NE_DRI_RDATA;
input  PLL0_NE_DRI_INTERRUPT;
output [10:0] PLL1_NE_DRI_CTRL;
input  [32:0] PLL1_NE_DRI_RDATA;
input  PLL1_NE_DRI_INTERRUPT;
output [10:0] PLL0_SE_DRI_CTRL;
input  [32:0] PLL0_SE_DRI_RDATA;
input  PLL0_SE_DRI_INTERRUPT;
output [10:0] PLL1_SE_DRI_CTRL;
input  [32:0] PLL1_SE_DRI_RDATA;
input  PLL1_SE_DRI_INTERRUPT;
output [10:0] PLL0_SW_DRI_CTRL;
input  [32:0] PLL0_SW_DRI_RDATA;
input  PLL0_SW_DRI_INTERRUPT;
output [10:0] PLL1_SW_DRI_CTRL;
input  [32:0] PLL1_SW_DRI_RDATA;
input  PLL1_SW_DRI_INTERRUPT;
output [10:0] DLL0_NW_DRI_CTRL;
input  [32:0] DLL0_NW_DRI_RDATA;
input  DLL0_NW_DRI_INTERRUPT;
output [10:0] DLL1_NW_DRI_CTRL;
input  [32:0] DLL1_NW_DRI_RDATA;
input  DLL1_NW_DRI_INTERRUPT;
output [10:0] DLL0_NE_DRI_CTRL;
input  [32:0] DLL0_NE_DRI_RDATA;
input  DLL0_NE_DRI_INTERRUPT;
output [10:0] DLL1_NE_DRI_CTRL;
input  [32:0] DLL1_NE_DRI_RDATA;
input  DLL1_NE_DRI_INTERRUPT;
output [10:0] DLL0_SE_DRI_CTRL;
input  [32:0] DLL0_SE_DRI_RDATA;
input  DLL0_SE_DRI_INTERRUPT;
output [10:0] DLL1_SE_DRI_CTRL;
input  [32:0] DLL1_SE_DRI_RDATA;
input  DLL1_SE_DRI_INTERRUPT;
output [10:0] DLL0_SW_DRI_CTRL;
input  [32:0] DLL0_SW_DRI_RDATA;
input  DLL0_SW_DRI_INTERRUPT;
output [10:0] DLL1_SW_DRI_CTRL;
input  [32:0] DLL1_SW_DRI_RDATA;
input  DLL1_SW_DRI_INTERRUPT;
output [10:0] CRYPTO_DRI_CTRL;
input  [32:0] CRYPTO_DRI_RDATA;
input  CRYPTO_DRI_INTERRUPT;
output DRI_CLK;
output [32:0] DRI_WDATA;
output DRI_ARST_N;

    wire gnd_net;
    
    GND gnd_inst (.Y(gnd_net));
    DRI I_DRI (.PRDATA({PRDATA[31], PRDATA[30], PRDATA[29], PRDATA[28], 
        PRDATA[27], PRDATA[26], PRDATA[25], PRDATA[24], PRDATA[23], 
        PRDATA[22], PRDATA[21], PRDATA[20], PRDATA[19], PRDATA[18], 
        PRDATA[17], PRDATA[16], PRDATA[15], PRDATA[14], PRDATA[13], 
        PRDATA[12], PRDATA[11], PRDATA[10], PRDATA[9], PRDATA[8], 
        PRDATA[7], PRDATA[6], PRDATA[5], PRDATA[4], PRDATA[3], 
        PRDATA[2], PRDATA[1], PRDATA[0]}), .PREADY(PREADY), .PSLVERR(
        PSLVERR), .PINTERRUPT(PINTERRUPT), .PTIMEOUT(PTIMEOUT), 
        .BUSERROR(BUSERROR), .PCLK(PCLK), .PSEL(PSEL), .PENABLE(
        PENABLE), .PWRITE(PWRITE), .PADDR({PADDR[28], PADDR[27], 
        PADDR[26], PADDR[25], PADDR[24], PADDR[23], PADDR[22], 
        PADDR[21], PADDR[20], PADDR[19], PADDR[18], PADDR[17], 
        PADDR[16], PADDR[15], PADDR[14], PADDR[13], PADDR[12], 
        PADDR[11], PADDR[10], PADDR[9], PADDR[8], PADDR[7], PADDR[6], 
        PADDR[5], PADDR[4], PADDR[3], PADDR[2], PADDR[1], PADDR[0]}), 
        .PSTRB({PSTRB[3], PSTRB[2], PSTRB[1], PSTRB[0]}), .PWDATA({
        PWDATA[31], PWDATA[30], PWDATA[29], PWDATA[28], PWDATA[27], 
        PWDATA[26], PWDATA[25], PWDATA[24], PWDATA[23], PWDATA[22], 
        PWDATA[21], PWDATA[20], PWDATA[19], PWDATA[18], PWDATA[17], 
        PWDATA[16], PWDATA[15], PWDATA[14], PWDATA[13], PWDATA[12], 
        PWDATA[11], PWDATA[10], PWDATA[9], PWDATA[8], PWDATA[7], 
        PWDATA[6], PWDATA[5], PWDATA[4], PWDATA[3], PWDATA[2], 
        PWDATA[1], PWDATA[0]}), .PRESETN(PRESETN), .DRI_CLK(DRI_CLK), 
        .DRI_WDATA({DRI_WDATA[32], DRI_WDATA[31], DRI_WDATA[30], 
        DRI_WDATA[29], DRI_WDATA[28], DRI_WDATA[27], DRI_WDATA[26], 
        DRI_WDATA[25], DRI_WDATA[24], DRI_WDATA[23], DRI_WDATA[22], 
        DRI_WDATA[21], DRI_WDATA[20], DRI_WDATA[19], DRI_WDATA[18], 
        DRI_WDATA[17], DRI_WDATA[16], DRI_WDATA[15], DRI_WDATA[14], 
        DRI_WDATA[13], DRI_WDATA[12], DRI_WDATA[11], DRI_WDATA[10], 
        DRI_WDATA[9], DRI_WDATA[8], DRI_WDATA[7], DRI_WDATA[6], 
        DRI_WDATA[5], DRI_WDATA[4], DRI_WDATA[3], DRI_WDATA[2], 
        DRI_WDATA[1], DRI_WDATA[0]}), .DRI_ARST_N(DRI_ARST_N), 
        .Q4_LANE0_DRI_CTRL({Q4_LANE0_DRI_CTRL[10], 
        Q4_LANE0_DRI_CTRL[9], Q4_LANE0_DRI_CTRL[8], 
        Q4_LANE0_DRI_CTRL[7], Q4_LANE0_DRI_CTRL[6], 
        Q4_LANE0_DRI_CTRL[5], Q4_LANE0_DRI_CTRL[4], 
        Q4_LANE0_DRI_CTRL[3], Q4_LANE0_DRI_CTRL[2], 
        Q4_LANE0_DRI_CTRL[1], Q4_LANE0_DRI_CTRL[0]}), 
        .Q4_LANE0_DRI_RDATA({Q4_LANE0_DRI_RDATA[32], 
        Q4_LANE0_DRI_RDATA[31], Q4_LANE0_DRI_RDATA[30], 
        Q4_LANE0_DRI_RDATA[29], Q4_LANE0_DRI_RDATA[28], 
        Q4_LANE0_DRI_RDATA[27], Q4_LANE0_DRI_RDATA[26], 
        Q4_LANE0_DRI_RDATA[25], Q4_LANE0_DRI_RDATA[24], 
        Q4_LANE0_DRI_RDATA[23], Q4_LANE0_DRI_RDATA[22], 
        Q4_LANE0_DRI_RDATA[21], Q4_LANE0_DRI_RDATA[20], 
        Q4_LANE0_DRI_RDATA[19], Q4_LANE0_DRI_RDATA[18], 
        Q4_LANE0_DRI_RDATA[17], Q4_LANE0_DRI_RDATA[16], 
        Q4_LANE0_DRI_RDATA[15], Q4_LANE0_DRI_RDATA[14], 
        Q4_LANE0_DRI_RDATA[13], Q4_LANE0_DRI_RDATA[12], 
        Q4_LANE0_DRI_RDATA[11], Q4_LANE0_DRI_RDATA[10], 
        Q4_LANE0_DRI_RDATA[9], Q4_LANE0_DRI_RDATA[8], 
        Q4_LANE0_DRI_RDATA[7], Q4_LANE0_DRI_RDATA[6], 
        Q4_LANE0_DRI_RDATA[5], Q4_LANE0_DRI_RDATA[4], 
        Q4_LANE0_DRI_RDATA[3], Q4_LANE0_DRI_RDATA[2], 
        Q4_LANE0_DRI_RDATA[1], Q4_LANE0_DRI_RDATA[0]}), 
        .Q4_LANE0_DRI_INTERRUPT(Q4_LANE0_DRI_INTERRUPT), 
        .Q4_LANE1_DRI_CTRL({Q4_LANE1_DRI_CTRL[10], 
        Q4_LANE1_DRI_CTRL[9], Q4_LANE1_DRI_CTRL[8], 
        Q4_LANE1_DRI_CTRL[7], Q4_LANE1_DRI_CTRL[6], 
        Q4_LANE1_DRI_CTRL[5], Q4_LANE1_DRI_CTRL[4], 
        Q4_LANE1_DRI_CTRL[3], Q4_LANE1_DRI_CTRL[2], 
        Q4_LANE1_DRI_CTRL[1], Q4_LANE1_DRI_CTRL[0]}), 
        .Q4_LANE1_DRI_RDATA({Q4_LANE1_DRI_RDATA[32], 
        Q4_LANE1_DRI_RDATA[31], Q4_LANE1_DRI_RDATA[30], 
        Q4_LANE1_DRI_RDATA[29], Q4_LANE1_DRI_RDATA[28], 
        Q4_LANE1_DRI_RDATA[27], Q4_LANE1_DRI_RDATA[26], 
        Q4_LANE1_DRI_RDATA[25], Q4_LANE1_DRI_RDATA[24], 
        Q4_LANE1_DRI_RDATA[23], Q4_LANE1_DRI_RDATA[22], 
        Q4_LANE1_DRI_RDATA[21], Q4_LANE1_DRI_RDATA[20], 
        Q4_LANE1_DRI_RDATA[19], Q4_LANE1_DRI_RDATA[18], 
        Q4_LANE1_DRI_RDATA[17], Q4_LANE1_DRI_RDATA[16], 
        Q4_LANE1_DRI_RDATA[15], Q4_LANE1_DRI_RDATA[14], 
        Q4_LANE1_DRI_RDATA[13], Q4_LANE1_DRI_RDATA[12], 
        Q4_LANE1_DRI_RDATA[11], Q4_LANE1_DRI_RDATA[10], 
        Q4_LANE1_DRI_RDATA[9], Q4_LANE1_DRI_RDATA[8], 
        Q4_LANE1_DRI_RDATA[7], Q4_LANE1_DRI_RDATA[6], 
        Q4_LANE1_DRI_RDATA[5], Q4_LANE1_DRI_RDATA[4], 
        Q4_LANE1_DRI_RDATA[3], Q4_LANE1_DRI_RDATA[2], 
        Q4_LANE1_DRI_RDATA[1], Q4_LANE1_DRI_RDATA[0]}), 
        .Q4_LANE1_DRI_INTERRUPT(Q4_LANE1_DRI_INTERRUPT), 
        .Q4_LANE2_DRI_CTRL({Q4_LANE2_DRI_CTRL[10], 
        Q4_LANE2_DRI_CTRL[9], Q4_LANE2_DRI_CTRL[8], 
        Q4_LANE2_DRI_CTRL[7], Q4_LANE2_DRI_CTRL[6], 
        Q4_LANE2_DRI_CTRL[5], Q4_LANE2_DRI_CTRL[4], 
        Q4_LANE2_DRI_CTRL[3], Q4_LANE2_DRI_CTRL[2], 
        Q4_LANE2_DRI_CTRL[1], Q4_LANE2_DRI_CTRL[0]}), 
        .Q4_LANE2_DRI_RDATA({Q4_LANE2_DRI_RDATA[32], 
        Q4_LANE2_DRI_RDATA[31], Q4_LANE2_DRI_RDATA[30], 
        Q4_LANE2_DRI_RDATA[29], Q4_LANE2_DRI_RDATA[28], 
        Q4_LANE2_DRI_RDATA[27], Q4_LANE2_DRI_RDATA[26], 
        Q4_LANE2_DRI_RDATA[25], Q4_LANE2_DRI_RDATA[24], 
        Q4_LANE2_DRI_RDATA[23], Q4_LANE2_DRI_RDATA[22], 
        Q4_LANE2_DRI_RDATA[21], Q4_LANE2_DRI_RDATA[20], 
        Q4_LANE2_DRI_RDATA[19], Q4_LANE2_DRI_RDATA[18], 
        Q4_LANE2_DRI_RDATA[17], Q4_LANE2_DRI_RDATA[16], 
        Q4_LANE2_DRI_RDATA[15], Q4_LANE2_DRI_RDATA[14], 
        Q4_LANE2_DRI_RDATA[13], Q4_LANE2_DRI_RDATA[12], 
        Q4_LANE2_DRI_RDATA[11], Q4_LANE2_DRI_RDATA[10], 
        Q4_LANE2_DRI_RDATA[9], Q4_LANE2_DRI_RDATA[8], 
        Q4_LANE2_DRI_RDATA[7], Q4_LANE2_DRI_RDATA[6], 
        Q4_LANE2_DRI_RDATA[5], Q4_LANE2_DRI_RDATA[4], 
        Q4_LANE2_DRI_RDATA[3], Q4_LANE2_DRI_RDATA[2], 
        Q4_LANE2_DRI_RDATA[1], Q4_LANE2_DRI_RDATA[0]}), 
        .Q4_LANE2_DRI_INTERRUPT(Q4_LANE2_DRI_INTERRUPT), 
        .Q4_LANE3_DRI_CTRL({Q4_LANE3_DRI_CTRL[10], 
        Q4_LANE3_DRI_CTRL[9], Q4_LANE3_DRI_CTRL[8], 
        Q4_LANE3_DRI_CTRL[7], Q4_LANE3_DRI_CTRL[6], 
        Q4_LANE3_DRI_CTRL[5], Q4_LANE3_DRI_CTRL[4], 
        Q4_LANE3_DRI_CTRL[3], Q4_LANE3_DRI_CTRL[2], 
        Q4_LANE3_DRI_CTRL[1], Q4_LANE3_DRI_CTRL[0]}), 
        .Q4_LANE3_DRI_RDATA({Q4_LANE3_DRI_RDATA[32], 
        Q4_LANE3_DRI_RDATA[31], Q4_LANE3_DRI_RDATA[30], 
        Q4_LANE3_DRI_RDATA[29], Q4_LANE3_DRI_RDATA[28], 
        Q4_LANE3_DRI_RDATA[27], Q4_LANE3_DRI_RDATA[26], 
        Q4_LANE3_DRI_RDATA[25], Q4_LANE3_DRI_RDATA[24], 
        Q4_LANE3_DRI_RDATA[23], Q4_LANE3_DRI_RDATA[22], 
        Q4_LANE3_DRI_RDATA[21], Q4_LANE3_DRI_RDATA[20], 
        Q4_LANE3_DRI_RDATA[19], Q4_LANE3_DRI_RDATA[18], 
        Q4_LANE3_DRI_RDATA[17], Q4_LANE3_DRI_RDATA[16], 
        Q4_LANE3_DRI_RDATA[15], Q4_LANE3_DRI_RDATA[14], 
        Q4_LANE3_DRI_RDATA[13], Q4_LANE3_DRI_RDATA[12], 
        Q4_LANE3_DRI_RDATA[11], Q4_LANE3_DRI_RDATA[10], 
        Q4_LANE3_DRI_RDATA[9], Q4_LANE3_DRI_RDATA[8], 
        Q4_LANE3_DRI_RDATA[7], Q4_LANE3_DRI_RDATA[6], 
        Q4_LANE3_DRI_RDATA[5], Q4_LANE3_DRI_RDATA[4], 
        Q4_LANE3_DRI_RDATA[3], Q4_LANE3_DRI_RDATA[2], 
        Q4_LANE3_DRI_RDATA[1], Q4_LANE3_DRI_RDATA[0]}), 
        .Q4_LANE3_DRI_INTERRUPT(Q4_LANE3_DRI_INTERRUPT), 
        .Q2_LANE0_DRI_CTRL({Q2_LANE0_DRI_CTRL[10], 
        Q2_LANE0_DRI_CTRL[9], Q2_LANE0_DRI_CTRL[8], 
        Q2_LANE0_DRI_CTRL[7], Q2_LANE0_DRI_CTRL[6], 
        Q2_LANE0_DRI_CTRL[5], Q2_LANE0_DRI_CTRL[4], 
        Q2_LANE0_DRI_CTRL[3], Q2_LANE0_DRI_CTRL[2], 
        Q2_LANE0_DRI_CTRL[1], Q2_LANE0_DRI_CTRL[0]}), 
        .Q2_LANE0_DRI_RDATA({Q2_LANE0_DRI_RDATA[32], 
        Q2_LANE0_DRI_RDATA[31], Q2_LANE0_DRI_RDATA[30], 
        Q2_LANE0_DRI_RDATA[29], Q2_LANE0_DRI_RDATA[28], 
        Q2_LANE0_DRI_RDATA[27], Q2_LANE0_DRI_RDATA[26], 
        Q2_LANE0_DRI_RDATA[25], Q2_LANE0_DRI_RDATA[24], 
        Q2_LANE0_DRI_RDATA[23], Q2_LANE0_DRI_RDATA[22], 
        Q2_LANE0_DRI_RDATA[21], Q2_LANE0_DRI_RDATA[20], 
        Q2_LANE0_DRI_RDATA[19], Q2_LANE0_DRI_RDATA[18], 
        Q2_LANE0_DRI_RDATA[17], Q2_LANE0_DRI_RDATA[16], 
        Q2_LANE0_DRI_RDATA[15], Q2_LANE0_DRI_RDATA[14], 
        Q2_LANE0_DRI_RDATA[13], Q2_LANE0_DRI_RDATA[12], 
        Q2_LANE0_DRI_RDATA[11], Q2_LANE0_DRI_RDATA[10], 
        Q2_LANE0_DRI_RDATA[9], Q2_LANE0_DRI_RDATA[8], 
        Q2_LANE0_DRI_RDATA[7], Q2_LANE0_DRI_RDATA[6], 
        Q2_LANE0_DRI_RDATA[5], Q2_LANE0_DRI_RDATA[4], 
        Q2_LANE0_DRI_RDATA[3], Q2_LANE0_DRI_RDATA[2], 
        Q2_LANE0_DRI_RDATA[1], Q2_LANE0_DRI_RDATA[0]}), 
        .Q2_LANE0_DRI_INTERRUPT(Q2_LANE0_DRI_INTERRUPT), 
        .Q2_LANE1_DRI_CTRL({Q2_LANE1_DRI_CTRL[10], 
        Q2_LANE1_DRI_CTRL[9], Q2_LANE1_DRI_CTRL[8], 
        Q2_LANE1_DRI_CTRL[7], Q2_LANE1_DRI_CTRL[6], 
        Q2_LANE1_DRI_CTRL[5], Q2_LANE1_DRI_CTRL[4], 
        Q2_LANE1_DRI_CTRL[3], Q2_LANE1_DRI_CTRL[2], 
        Q2_LANE1_DRI_CTRL[1], Q2_LANE1_DRI_CTRL[0]}), 
        .Q2_LANE1_DRI_RDATA({Q2_LANE1_DRI_RDATA[32], 
        Q2_LANE1_DRI_RDATA[31], Q2_LANE1_DRI_RDATA[30], 
        Q2_LANE1_DRI_RDATA[29], Q2_LANE1_DRI_RDATA[28], 
        Q2_LANE1_DRI_RDATA[27], Q2_LANE1_DRI_RDATA[26], 
        Q2_LANE1_DRI_RDATA[25], Q2_LANE1_DRI_RDATA[24], 
        Q2_LANE1_DRI_RDATA[23], Q2_LANE1_DRI_RDATA[22], 
        Q2_LANE1_DRI_RDATA[21], Q2_LANE1_DRI_RDATA[20], 
        Q2_LANE1_DRI_RDATA[19], Q2_LANE1_DRI_RDATA[18], 
        Q2_LANE1_DRI_RDATA[17], Q2_LANE1_DRI_RDATA[16], 
        Q2_LANE1_DRI_RDATA[15], Q2_LANE1_DRI_RDATA[14], 
        Q2_LANE1_DRI_RDATA[13], Q2_LANE1_DRI_RDATA[12], 
        Q2_LANE1_DRI_RDATA[11], Q2_LANE1_DRI_RDATA[10], 
        Q2_LANE1_DRI_RDATA[9], Q2_LANE1_DRI_RDATA[8], 
        Q2_LANE1_DRI_RDATA[7], Q2_LANE1_DRI_RDATA[6], 
        Q2_LANE1_DRI_RDATA[5], Q2_LANE1_DRI_RDATA[4], 
        Q2_LANE1_DRI_RDATA[3], Q2_LANE1_DRI_RDATA[2], 
        Q2_LANE1_DRI_RDATA[1], Q2_LANE1_DRI_RDATA[0]}), 
        .Q2_LANE1_DRI_INTERRUPT(Q2_LANE1_DRI_INTERRUPT), 
        .Q2_LANE2_DRI_CTRL({Q2_LANE2_DRI_CTRL[10], 
        Q2_LANE2_DRI_CTRL[9], Q2_LANE2_DRI_CTRL[8], 
        Q2_LANE2_DRI_CTRL[7], Q2_LANE2_DRI_CTRL[6], 
        Q2_LANE2_DRI_CTRL[5], Q2_LANE2_DRI_CTRL[4], 
        Q2_LANE2_DRI_CTRL[3], Q2_LANE2_DRI_CTRL[2], 
        Q2_LANE2_DRI_CTRL[1], Q2_LANE2_DRI_CTRL[0]}), 
        .Q2_LANE2_DRI_RDATA({Q2_LANE2_DRI_RDATA[32], 
        Q2_LANE2_DRI_RDATA[31], Q2_LANE2_DRI_RDATA[30], 
        Q2_LANE2_DRI_RDATA[29], Q2_LANE2_DRI_RDATA[28], 
        Q2_LANE2_DRI_RDATA[27], Q2_LANE2_DRI_RDATA[26], 
        Q2_LANE2_DRI_RDATA[25], Q2_LANE2_DRI_RDATA[24], 
        Q2_LANE2_DRI_RDATA[23], Q2_LANE2_DRI_RDATA[22], 
        Q2_LANE2_DRI_RDATA[21], Q2_LANE2_DRI_RDATA[20], 
        Q2_LANE2_DRI_RDATA[19], Q2_LANE2_DRI_RDATA[18], 
        Q2_LANE2_DRI_RDATA[17], Q2_LANE2_DRI_RDATA[16], 
        Q2_LANE2_DRI_RDATA[15], Q2_LANE2_DRI_RDATA[14], 
        Q2_LANE2_DRI_RDATA[13], Q2_LANE2_DRI_RDATA[12], 
        Q2_LANE2_DRI_RDATA[11], Q2_LANE2_DRI_RDATA[10], 
        Q2_LANE2_DRI_RDATA[9], Q2_LANE2_DRI_RDATA[8], 
        Q2_LANE2_DRI_RDATA[7], Q2_LANE2_DRI_RDATA[6], 
        Q2_LANE2_DRI_RDATA[5], Q2_LANE2_DRI_RDATA[4], 
        Q2_LANE2_DRI_RDATA[3], Q2_LANE2_DRI_RDATA[2], 
        Q2_LANE2_DRI_RDATA[1], Q2_LANE2_DRI_RDATA[0]}), 
        .Q2_LANE2_DRI_INTERRUPT(Q2_LANE2_DRI_INTERRUPT), 
        .Q2_LANE3_DRI_CTRL({Q2_LANE3_DRI_CTRL[10], 
        Q2_LANE3_DRI_CTRL[9], Q2_LANE3_DRI_CTRL[8], 
        Q2_LANE3_DRI_CTRL[7], Q2_LANE3_DRI_CTRL[6], 
        Q2_LANE3_DRI_CTRL[5], Q2_LANE3_DRI_CTRL[4], 
        Q2_LANE3_DRI_CTRL[3], Q2_LANE3_DRI_CTRL[2], 
        Q2_LANE3_DRI_CTRL[1], Q2_LANE3_DRI_CTRL[0]}), 
        .Q2_LANE3_DRI_RDATA({Q2_LANE3_DRI_RDATA[32], 
        Q2_LANE3_DRI_RDATA[31], Q2_LANE3_DRI_RDATA[30], 
        Q2_LANE3_DRI_RDATA[29], Q2_LANE3_DRI_RDATA[28], 
        Q2_LANE3_DRI_RDATA[27], Q2_LANE3_DRI_RDATA[26], 
        Q2_LANE3_DRI_RDATA[25], Q2_LANE3_DRI_RDATA[24], 
        Q2_LANE3_DRI_RDATA[23], Q2_LANE3_DRI_RDATA[22], 
        Q2_LANE3_DRI_RDATA[21], Q2_LANE3_DRI_RDATA[20], 
        Q2_LANE3_DRI_RDATA[19], Q2_LANE3_DRI_RDATA[18], 
        Q2_LANE3_DRI_RDATA[17], Q2_LANE3_DRI_RDATA[16], 
        Q2_LANE3_DRI_RDATA[15], Q2_LANE3_DRI_RDATA[14], 
        Q2_LANE3_DRI_RDATA[13], Q2_LANE3_DRI_RDATA[12], 
        Q2_LANE3_DRI_RDATA[11], Q2_LANE3_DRI_RDATA[10], 
        Q2_LANE3_DRI_RDATA[9], Q2_LANE3_DRI_RDATA[8], 
        Q2_LANE3_DRI_RDATA[7], Q2_LANE3_DRI_RDATA[6], 
        Q2_LANE3_DRI_RDATA[5], Q2_LANE3_DRI_RDATA[4], 
        Q2_LANE3_DRI_RDATA[3], Q2_LANE3_DRI_RDATA[2], 
        Q2_LANE3_DRI_RDATA[1], Q2_LANE3_DRI_RDATA[0]}), 
        .Q2_LANE3_DRI_INTERRUPT(Q2_LANE3_DRI_INTERRUPT), 
        .Q0_LANE0_DRI_CTRL({Q0_LANE0_DRI_CTRL[10], 
        Q0_LANE0_DRI_CTRL[9], Q0_LANE0_DRI_CTRL[8], 
        Q0_LANE0_DRI_CTRL[7], Q0_LANE0_DRI_CTRL[6], 
        Q0_LANE0_DRI_CTRL[5], Q0_LANE0_DRI_CTRL[4], 
        Q0_LANE0_DRI_CTRL[3], Q0_LANE0_DRI_CTRL[2], 
        Q0_LANE0_DRI_CTRL[1], Q0_LANE0_DRI_CTRL[0]}), 
        .Q0_LANE0_DRI_RDATA({Q0_LANE0_DRI_RDATA[32], 
        Q0_LANE0_DRI_RDATA[31], Q0_LANE0_DRI_RDATA[30], 
        Q0_LANE0_DRI_RDATA[29], Q0_LANE0_DRI_RDATA[28], 
        Q0_LANE0_DRI_RDATA[27], Q0_LANE0_DRI_RDATA[26], 
        Q0_LANE0_DRI_RDATA[25], Q0_LANE0_DRI_RDATA[24], 
        Q0_LANE0_DRI_RDATA[23], Q0_LANE0_DRI_RDATA[22], 
        Q0_LANE0_DRI_RDATA[21], Q0_LANE0_DRI_RDATA[20], 
        Q0_LANE0_DRI_RDATA[19], Q0_LANE0_DRI_RDATA[18], 
        Q0_LANE0_DRI_RDATA[17], Q0_LANE0_DRI_RDATA[16], 
        Q0_LANE0_DRI_RDATA[15], Q0_LANE0_DRI_RDATA[14], 
        Q0_LANE0_DRI_RDATA[13], Q0_LANE0_DRI_RDATA[12], 
        Q0_LANE0_DRI_RDATA[11], Q0_LANE0_DRI_RDATA[10], 
        Q0_LANE0_DRI_RDATA[9], Q0_LANE0_DRI_RDATA[8], 
        Q0_LANE0_DRI_RDATA[7], Q0_LANE0_DRI_RDATA[6], 
        Q0_LANE0_DRI_RDATA[5], Q0_LANE0_DRI_RDATA[4], 
        Q0_LANE0_DRI_RDATA[3], Q0_LANE0_DRI_RDATA[2], 
        Q0_LANE0_DRI_RDATA[1], Q0_LANE0_DRI_RDATA[0]}), 
        .Q0_LANE0_DRI_INTERRUPT(Q0_LANE0_DRI_INTERRUPT), 
        .Q0_LANE1_DRI_CTRL({Q0_LANE1_DRI_CTRL[10], 
        Q0_LANE1_DRI_CTRL[9], Q0_LANE1_DRI_CTRL[8], 
        Q0_LANE1_DRI_CTRL[7], Q0_LANE1_DRI_CTRL[6], 
        Q0_LANE1_DRI_CTRL[5], Q0_LANE1_DRI_CTRL[4], 
        Q0_LANE1_DRI_CTRL[3], Q0_LANE1_DRI_CTRL[2], 
        Q0_LANE1_DRI_CTRL[1], Q0_LANE1_DRI_CTRL[0]}), 
        .Q0_LANE1_DRI_RDATA({Q0_LANE1_DRI_RDATA[32], 
        Q0_LANE1_DRI_RDATA[31], Q0_LANE1_DRI_RDATA[30], 
        Q0_LANE1_DRI_RDATA[29], Q0_LANE1_DRI_RDATA[28], 
        Q0_LANE1_DRI_RDATA[27], Q0_LANE1_DRI_RDATA[26], 
        Q0_LANE1_DRI_RDATA[25], Q0_LANE1_DRI_RDATA[24], 
        Q0_LANE1_DRI_RDATA[23], Q0_LANE1_DRI_RDATA[22], 
        Q0_LANE1_DRI_RDATA[21], Q0_LANE1_DRI_RDATA[20], 
        Q0_LANE1_DRI_RDATA[19], Q0_LANE1_DRI_RDATA[18], 
        Q0_LANE1_DRI_RDATA[17], Q0_LANE1_DRI_RDATA[16], 
        Q0_LANE1_DRI_RDATA[15], Q0_LANE1_DRI_RDATA[14], 
        Q0_LANE1_DRI_RDATA[13], Q0_LANE1_DRI_RDATA[12], 
        Q0_LANE1_DRI_RDATA[11], Q0_LANE1_DRI_RDATA[10], 
        Q0_LANE1_DRI_RDATA[9], Q0_LANE1_DRI_RDATA[8], 
        Q0_LANE1_DRI_RDATA[7], Q0_LANE1_DRI_RDATA[6], 
        Q0_LANE1_DRI_RDATA[5], Q0_LANE1_DRI_RDATA[4], 
        Q0_LANE1_DRI_RDATA[3], Q0_LANE1_DRI_RDATA[2], 
        Q0_LANE1_DRI_RDATA[1], Q0_LANE1_DRI_RDATA[0]}), 
        .Q0_LANE1_DRI_INTERRUPT(Q0_LANE1_DRI_INTERRUPT), 
        .Q0_LANE2_DRI_CTRL({Q0_LANE2_DRI_CTRL[10], 
        Q0_LANE2_DRI_CTRL[9], Q0_LANE2_DRI_CTRL[8], 
        Q0_LANE2_DRI_CTRL[7], Q0_LANE2_DRI_CTRL[6], 
        Q0_LANE2_DRI_CTRL[5], Q0_LANE2_DRI_CTRL[4], 
        Q0_LANE2_DRI_CTRL[3], Q0_LANE2_DRI_CTRL[2], 
        Q0_LANE2_DRI_CTRL[1], Q0_LANE2_DRI_CTRL[0]}), 
        .Q0_LANE2_DRI_RDATA({Q0_LANE2_DRI_RDATA[32], 
        Q0_LANE2_DRI_RDATA[31], Q0_LANE2_DRI_RDATA[30], 
        Q0_LANE2_DRI_RDATA[29], Q0_LANE2_DRI_RDATA[28], 
        Q0_LANE2_DRI_RDATA[27], Q0_LANE2_DRI_RDATA[26], 
        Q0_LANE2_DRI_RDATA[25], Q0_LANE2_DRI_RDATA[24], 
        Q0_LANE2_DRI_RDATA[23], Q0_LANE2_DRI_RDATA[22], 
        Q0_LANE2_DRI_RDATA[21], Q0_LANE2_DRI_RDATA[20], 
        Q0_LANE2_DRI_RDATA[19], Q0_LANE2_DRI_RDATA[18], 
        Q0_LANE2_DRI_RDATA[17], Q0_LANE2_DRI_RDATA[16], 
        Q0_LANE2_DRI_RDATA[15], Q0_LANE2_DRI_RDATA[14], 
        Q0_LANE2_DRI_RDATA[13], Q0_LANE2_DRI_RDATA[12], 
        Q0_LANE2_DRI_RDATA[11], Q0_LANE2_DRI_RDATA[10], 
        Q0_LANE2_DRI_RDATA[9], Q0_LANE2_DRI_RDATA[8], 
        Q0_LANE2_DRI_RDATA[7], Q0_LANE2_DRI_RDATA[6], 
        Q0_LANE2_DRI_RDATA[5], Q0_LANE2_DRI_RDATA[4], 
        Q0_LANE2_DRI_RDATA[3], Q0_LANE2_DRI_RDATA[2], 
        Q0_LANE2_DRI_RDATA[1], Q0_LANE2_DRI_RDATA[0]}), 
        .Q0_LANE2_DRI_INTERRUPT(Q0_LANE2_DRI_INTERRUPT), 
        .Q0_LANE3_DRI_CTRL({Q0_LANE3_DRI_CTRL[10], 
        Q0_LANE3_DRI_CTRL[9], Q0_LANE3_DRI_CTRL[8], 
        Q0_LANE3_DRI_CTRL[7], Q0_LANE3_DRI_CTRL[6], 
        Q0_LANE3_DRI_CTRL[5], Q0_LANE3_DRI_CTRL[4], 
        Q0_LANE3_DRI_CTRL[3], Q0_LANE3_DRI_CTRL[2], 
        Q0_LANE3_DRI_CTRL[1], Q0_LANE3_DRI_CTRL[0]}), 
        .Q0_LANE3_DRI_RDATA({Q0_LANE3_DRI_RDATA[32], 
        Q0_LANE3_DRI_RDATA[31], Q0_LANE3_DRI_RDATA[30], 
        Q0_LANE3_DRI_RDATA[29], Q0_LANE3_DRI_RDATA[28], 
        Q0_LANE3_DRI_RDATA[27], Q0_LANE3_DRI_RDATA[26], 
        Q0_LANE3_DRI_RDATA[25], Q0_LANE3_DRI_RDATA[24], 
        Q0_LANE3_DRI_RDATA[23], Q0_LANE3_DRI_RDATA[22], 
        Q0_LANE3_DRI_RDATA[21], Q0_LANE3_DRI_RDATA[20], 
        Q0_LANE3_DRI_RDATA[19], Q0_LANE3_DRI_RDATA[18], 
        Q0_LANE3_DRI_RDATA[17], Q0_LANE3_DRI_RDATA[16], 
        Q0_LANE3_DRI_RDATA[15], Q0_LANE3_DRI_RDATA[14], 
        Q0_LANE3_DRI_RDATA[13], Q0_LANE3_DRI_RDATA[12], 
        Q0_LANE3_DRI_RDATA[11], Q0_LANE3_DRI_RDATA[10], 
        Q0_LANE3_DRI_RDATA[9], Q0_LANE3_DRI_RDATA[8], 
        Q0_LANE3_DRI_RDATA[7], Q0_LANE3_DRI_RDATA[6], 
        Q0_LANE3_DRI_RDATA[5], Q0_LANE3_DRI_RDATA[4], 
        Q0_LANE3_DRI_RDATA[3], Q0_LANE3_DRI_RDATA[2], 
        Q0_LANE3_DRI_RDATA[1], Q0_LANE3_DRI_RDATA[0]}), 
        .Q0_LANE3_DRI_INTERRUPT(Q0_LANE3_DRI_INTERRUPT), 
        .Q1_LANE0_DRI_CTRL({Q1_LANE0_DRI_CTRL[10], 
        Q1_LANE0_DRI_CTRL[9], Q1_LANE0_DRI_CTRL[8], 
        Q1_LANE0_DRI_CTRL[7], Q1_LANE0_DRI_CTRL[6], 
        Q1_LANE0_DRI_CTRL[5], Q1_LANE0_DRI_CTRL[4], 
        Q1_LANE0_DRI_CTRL[3], Q1_LANE0_DRI_CTRL[2], 
        Q1_LANE0_DRI_CTRL[1], Q1_LANE0_DRI_CTRL[0]}), 
        .Q1_LANE0_DRI_RDATA({Q1_LANE0_DRI_RDATA[32], 
        Q1_LANE0_DRI_RDATA[31], Q1_LANE0_DRI_RDATA[30], 
        Q1_LANE0_DRI_RDATA[29], Q1_LANE0_DRI_RDATA[28], 
        Q1_LANE0_DRI_RDATA[27], Q1_LANE0_DRI_RDATA[26], 
        Q1_LANE0_DRI_RDATA[25], Q1_LANE0_DRI_RDATA[24], 
        Q1_LANE0_DRI_RDATA[23], Q1_LANE0_DRI_RDATA[22], 
        Q1_LANE0_DRI_RDATA[21], Q1_LANE0_DRI_RDATA[20], 
        Q1_LANE0_DRI_RDATA[19], Q1_LANE0_DRI_RDATA[18], 
        Q1_LANE0_DRI_RDATA[17], Q1_LANE0_DRI_RDATA[16], 
        Q1_LANE0_DRI_RDATA[15], Q1_LANE0_DRI_RDATA[14], 
        Q1_LANE0_DRI_RDATA[13], Q1_LANE0_DRI_RDATA[12], 
        Q1_LANE0_DRI_RDATA[11], Q1_LANE0_DRI_RDATA[10], 
        Q1_LANE0_DRI_RDATA[9], Q1_LANE0_DRI_RDATA[8], 
        Q1_LANE0_DRI_RDATA[7], Q1_LANE0_DRI_RDATA[6], 
        Q1_LANE0_DRI_RDATA[5], Q1_LANE0_DRI_RDATA[4], 
        Q1_LANE0_DRI_RDATA[3], Q1_LANE0_DRI_RDATA[2], 
        Q1_LANE0_DRI_RDATA[1], Q1_LANE0_DRI_RDATA[0]}), 
        .Q1_LANE0_DRI_INTERRUPT(Q1_LANE0_DRI_INTERRUPT), 
        .Q1_LANE1_DRI_CTRL({Q1_LANE1_DRI_CTRL[10], 
        Q1_LANE1_DRI_CTRL[9], Q1_LANE1_DRI_CTRL[8], 
        Q1_LANE1_DRI_CTRL[7], Q1_LANE1_DRI_CTRL[6], 
        Q1_LANE1_DRI_CTRL[5], Q1_LANE1_DRI_CTRL[4], 
        Q1_LANE1_DRI_CTRL[3], Q1_LANE1_DRI_CTRL[2], 
        Q1_LANE1_DRI_CTRL[1], Q1_LANE1_DRI_CTRL[0]}), 
        .Q1_LANE1_DRI_RDATA({Q1_LANE1_DRI_RDATA[32], 
        Q1_LANE1_DRI_RDATA[31], Q1_LANE1_DRI_RDATA[30], 
        Q1_LANE1_DRI_RDATA[29], Q1_LANE1_DRI_RDATA[28], 
        Q1_LANE1_DRI_RDATA[27], Q1_LANE1_DRI_RDATA[26], 
        Q1_LANE1_DRI_RDATA[25], Q1_LANE1_DRI_RDATA[24], 
        Q1_LANE1_DRI_RDATA[23], Q1_LANE1_DRI_RDATA[22], 
        Q1_LANE1_DRI_RDATA[21], Q1_LANE1_DRI_RDATA[20], 
        Q1_LANE1_DRI_RDATA[19], Q1_LANE1_DRI_RDATA[18], 
        Q1_LANE1_DRI_RDATA[17], Q1_LANE1_DRI_RDATA[16], 
        Q1_LANE1_DRI_RDATA[15], Q1_LANE1_DRI_RDATA[14], 
        Q1_LANE1_DRI_RDATA[13], Q1_LANE1_DRI_RDATA[12], 
        Q1_LANE1_DRI_RDATA[11], Q1_LANE1_DRI_RDATA[10], 
        Q1_LANE1_DRI_RDATA[9], Q1_LANE1_DRI_RDATA[8], 
        Q1_LANE1_DRI_RDATA[7], Q1_LANE1_DRI_RDATA[6], 
        Q1_LANE1_DRI_RDATA[5], Q1_LANE1_DRI_RDATA[4], 
        Q1_LANE1_DRI_RDATA[3], Q1_LANE1_DRI_RDATA[2], 
        Q1_LANE1_DRI_RDATA[1], Q1_LANE1_DRI_RDATA[0]}), 
        .Q1_LANE1_DRI_INTERRUPT(Q1_LANE1_DRI_INTERRUPT), 
        .Q1_LANE2_DRI_CTRL({Q1_LANE2_DRI_CTRL[10], 
        Q1_LANE2_DRI_CTRL[9], Q1_LANE2_DRI_CTRL[8], 
        Q1_LANE2_DRI_CTRL[7], Q1_LANE2_DRI_CTRL[6], 
        Q1_LANE2_DRI_CTRL[5], Q1_LANE2_DRI_CTRL[4], 
        Q1_LANE2_DRI_CTRL[3], Q1_LANE2_DRI_CTRL[2], 
        Q1_LANE2_DRI_CTRL[1], Q1_LANE2_DRI_CTRL[0]}), 
        .Q1_LANE2_DRI_RDATA({Q1_LANE2_DRI_RDATA[32], 
        Q1_LANE2_DRI_RDATA[31], Q1_LANE2_DRI_RDATA[30], 
        Q1_LANE2_DRI_RDATA[29], Q1_LANE2_DRI_RDATA[28], 
        Q1_LANE2_DRI_RDATA[27], Q1_LANE2_DRI_RDATA[26], 
        Q1_LANE2_DRI_RDATA[25], Q1_LANE2_DRI_RDATA[24], 
        Q1_LANE2_DRI_RDATA[23], Q1_LANE2_DRI_RDATA[22], 
        Q1_LANE2_DRI_RDATA[21], Q1_LANE2_DRI_RDATA[20], 
        Q1_LANE2_DRI_RDATA[19], Q1_LANE2_DRI_RDATA[18], 
        Q1_LANE2_DRI_RDATA[17], Q1_LANE2_DRI_RDATA[16], 
        Q1_LANE2_DRI_RDATA[15], Q1_LANE2_DRI_RDATA[14], 
        Q1_LANE2_DRI_RDATA[13], Q1_LANE2_DRI_RDATA[12], 
        Q1_LANE2_DRI_RDATA[11], Q1_LANE2_DRI_RDATA[10], 
        Q1_LANE2_DRI_RDATA[9], Q1_LANE2_DRI_RDATA[8], 
        Q1_LANE2_DRI_RDATA[7], Q1_LANE2_DRI_RDATA[6], 
        Q1_LANE2_DRI_RDATA[5], Q1_LANE2_DRI_RDATA[4], 
        Q1_LANE2_DRI_RDATA[3], Q1_LANE2_DRI_RDATA[2], 
        Q1_LANE2_DRI_RDATA[1], Q1_LANE2_DRI_RDATA[0]}), 
        .Q1_LANE2_DRI_INTERRUPT(Q1_LANE2_DRI_INTERRUPT), 
        .Q1_LANE3_DRI_CTRL({Q1_LANE3_DRI_CTRL[10], 
        Q1_LANE3_DRI_CTRL[9], Q1_LANE3_DRI_CTRL[8], 
        Q1_LANE3_DRI_CTRL[7], Q1_LANE3_DRI_CTRL[6], 
        Q1_LANE3_DRI_CTRL[5], Q1_LANE3_DRI_CTRL[4], 
        Q1_LANE3_DRI_CTRL[3], Q1_LANE3_DRI_CTRL[2], 
        Q1_LANE3_DRI_CTRL[1], Q1_LANE3_DRI_CTRL[0]}), 
        .Q1_LANE3_DRI_RDATA({Q1_LANE3_DRI_RDATA[32], 
        Q1_LANE3_DRI_RDATA[31], Q1_LANE3_DRI_RDATA[30], 
        Q1_LANE3_DRI_RDATA[29], Q1_LANE3_DRI_RDATA[28], 
        Q1_LANE3_DRI_RDATA[27], Q1_LANE3_DRI_RDATA[26], 
        Q1_LANE3_DRI_RDATA[25], Q1_LANE3_DRI_RDATA[24], 
        Q1_LANE3_DRI_RDATA[23], Q1_LANE3_DRI_RDATA[22], 
        Q1_LANE3_DRI_RDATA[21], Q1_LANE3_DRI_RDATA[20], 
        Q1_LANE3_DRI_RDATA[19], Q1_LANE3_DRI_RDATA[18], 
        Q1_LANE3_DRI_RDATA[17], Q1_LANE3_DRI_RDATA[16], 
        Q1_LANE3_DRI_RDATA[15], Q1_LANE3_DRI_RDATA[14], 
        Q1_LANE3_DRI_RDATA[13], Q1_LANE3_DRI_RDATA[12], 
        Q1_LANE3_DRI_RDATA[11], Q1_LANE3_DRI_RDATA[10], 
        Q1_LANE3_DRI_RDATA[9], Q1_LANE3_DRI_RDATA[8], 
        Q1_LANE3_DRI_RDATA[7], Q1_LANE3_DRI_RDATA[6], 
        Q1_LANE3_DRI_RDATA[5], Q1_LANE3_DRI_RDATA[4], 
        Q1_LANE3_DRI_RDATA[3], Q1_LANE3_DRI_RDATA[2], 
        Q1_LANE3_DRI_RDATA[1], Q1_LANE3_DRI_RDATA[0]}), 
        .Q1_LANE3_DRI_INTERRUPT(Q1_LANE3_DRI_INTERRUPT), 
        .Q3_LANE0_DRI_CTRL({Q3_LANE0_DRI_CTRL[10], 
        Q3_LANE0_DRI_CTRL[9], Q3_LANE0_DRI_CTRL[8], 
        Q3_LANE0_DRI_CTRL[7], Q3_LANE0_DRI_CTRL[6], 
        Q3_LANE0_DRI_CTRL[5], Q3_LANE0_DRI_CTRL[4], 
        Q3_LANE0_DRI_CTRL[3], Q3_LANE0_DRI_CTRL[2], 
        Q3_LANE0_DRI_CTRL[1], Q3_LANE0_DRI_CTRL[0]}), 
        .Q3_LANE0_DRI_RDATA({Q3_LANE0_DRI_RDATA[32], 
        Q3_LANE0_DRI_RDATA[31], Q3_LANE0_DRI_RDATA[30], 
        Q3_LANE0_DRI_RDATA[29], Q3_LANE0_DRI_RDATA[28], 
        Q3_LANE0_DRI_RDATA[27], Q3_LANE0_DRI_RDATA[26], 
        Q3_LANE0_DRI_RDATA[25], Q3_LANE0_DRI_RDATA[24], 
        Q3_LANE0_DRI_RDATA[23], Q3_LANE0_DRI_RDATA[22], 
        Q3_LANE0_DRI_RDATA[21], Q3_LANE0_DRI_RDATA[20], 
        Q3_LANE0_DRI_RDATA[19], Q3_LANE0_DRI_RDATA[18], 
        Q3_LANE0_DRI_RDATA[17], Q3_LANE0_DRI_RDATA[16], 
        Q3_LANE0_DRI_RDATA[15], Q3_LANE0_DRI_RDATA[14], 
        Q3_LANE0_DRI_RDATA[13], Q3_LANE0_DRI_RDATA[12], 
        Q3_LANE0_DRI_RDATA[11], Q3_LANE0_DRI_RDATA[10], 
        Q3_LANE0_DRI_RDATA[9], Q3_LANE0_DRI_RDATA[8], 
        Q3_LANE0_DRI_RDATA[7], Q3_LANE0_DRI_RDATA[6], 
        Q3_LANE0_DRI_RDATA[5], Q3_LANE0_DRI_RDATA[4], 
        Q3_LANE0_DRI_RDATA[3], Q3_LANE0_DRI_RDATA[2], 
        Q3_LANE0_DRI_RDATA[1], Q3_LANE0_DRI_RDATA[0]}), 
        .Q3_LANE0_DRI_INTERRUPT(Q3_LANE0_DRI_INTERRUPT), 
        .Q3_LANE1_DRI_CTRL({Q3_LANE1_DRI_CTRL[10], 
        Q3_LANE1_DRI_CTRL[9], Q3_LANE1_DRI_CTRL[8], 
        Q3_LANE1_DRI_CTRL[7], Q3_LANE1_DRI_CTRL[6], 
        Q3_LANE1_DRI_CTRL[5], Q3_LANE1_DRI_CTRL[4], 
        Q3_LANE1_DRI_CTRL[3], Q3_LANE1_DRI_CTRL[2], 
        Q3_LANE1_DRI_CTRL[1], Q3_LANE1_DRI_CTRL[0]}), 
        .Q3_LANE1_DRI_RDATA({Q3_LANE1_DRI_RDATA[32], 
        Q3_LANE1_DRI_RDATA[31], Q3_LANE1_DRI_RDATA[30], 
        Q3_LANE1_DRI_RDATA[29], Q3_LANE1_DRI_RDATA[28], 
        Q3_LANE1_DRI_RDATA[27], Q3_LANE1_DRI_RDATA[26], 
        Q3_LANE1_DRI_RDATA[25], Q3_LANE1_DRI_RDATA[24], 
        Q3_LANE1_DRI_RDATA[23], Q3_LANE1_DRI_RDATA[22], 
        Q3_LANE1_DRI_RDATA[21], Q3_LANE1_DRI_RDATA[20], 
        Q3_LANE1_DRI_RDATA[19], Q3_LANE1_DRI_RDATA[18], 
        Q3_LANE1_DRI_RDATA[17], Q3_LANE1_DRI_RDATA[16], 
        Q3_LANE1_DRI_RDATA[15], Q3_LANE1_DRI_RDATA[14], 
        Q3_LANE1_DRI_RDATA[13], Q3_LANE1_DRI_RDATA[12], 
        Q3_LANE1_DRI_RDATA[11], Q3_LANE1_DRI_RDATA[10], 
        Q3_LANE1_DRI_RDATA[9], Q3_LANE1_DRI_RDATA[8], 
        Q3_LANE1_DRI_RDATA[7], Q3_LANE1_DRI_RDATA[6], 
        Q3_LANE1_DRI_RDATA[5], Q3_LANE1_DRI_RDATA[4], 
        Q3_LANE1_DRI_RDATA[3], Q3_LANE1_DRI_RDATA[2], 
        Q3_LANE1_DRI_RDATA[1], Q3_LANE1_DRI_RDATA[0]}), 
        .Q3_LANE1_DRI_INTERRUPT(Q3_LANE1_DRI_INTERRUPT), 
        .Q3_LANE2_DRI_CTRL({Q3_LANE2_DRI_CTRL[10], 
        Q3_LANE2_DRI_CTRL[9], Q3_LANE2_DRI_CTRL[8], 
        Q3_LANE2_DRI_CTRL[7], Q3_LANE2_DRI_CTRL[6], 
        Q3_LANE2_DRI_CTRL[5], Q3_LANE2_DRI_CTRL[4], 
        Q3_LANE2_DRI_CTRL[3], Q3_LANE2_DRI_CTRL[2], 
        Q3_LANE2_DRI_CTRL[1], Q3_LANE2_DRI_CTRL[0]}), 
        .Q3_LANE2_DRI_RDATA({Q3_LANE2_DRI_RDATA[32], 
        Q3_LANE2_DRI_RDATA[31], Q3_LANE2_DRI_RDATA[30], 
        Q3_LANE2_DRI_RDATA[29], Q3_LANE2_DRI_RDATA[28], 
        Q3_LANE2_DRI_RDATA[27], Q3_LANE2_DRI_RDATA[26], 
        Q3_LANE2_DRI_RDATA[25], Q3_LANE2_DRI_RDATA[24], 
        Q3_LANE2_DRI_RDATA[23], Q3_LANE2_DRI_RDATA[22], 
        Q3_LANE2_DRI_RDATA[21], Q3_LANE2_DRI_RDATA[20], 
        Q3_LANE2_DRI_RDATA[19], Q3_LANE2_DRI_RDATA[18], 
        Q3_LANE2_DRI_RDATA[17], Q3_LANE2_DRI_RDATA[16], 
        Q3_LANE2_DRI_RDATA[15], Q3_LANE2_DRI_RDATA[14], 
        Q3_LANE2_DRI_RDATA[13], Q3_LANE2_DRI_RDATA[12], 
        Q3_LANE2_DRI_RDATA[11], Q3_LANE2_DRI_RDATA[10], 
        Q3_LANE2_DRI_RDATA[9], Q3_LANE2_DRI_RDATA[8], 
        Q3_LANE2_DRI_RDATA[7], Q3_LANE2_DRI_RDATA[6], 
        Q3_LANE2_DRI_RDATA[5], Q3_LANE2_DRI_RDATA[4], 
        Q3_LANE2_DRI_RDATA[3], Q3_LANE2_DRI_RDATA[2], 
        Q3_LANE2_DRI_RDATA[1], Q3_LANE2_DRI_RDATA[0]}), 
        .Q3_LANE2_DRI_INTERRUPT(Q3_LANE2_DRI_INTERRUPT), 
        .Q3_LANE3_DRI_CTRL({Q3_LANE3_DRI_CTRL[10], 
        Q3_LANE3_DRI_CTRL[9], Q3_LANE3_DRI_CTRL[8], 
        Q3_LANE3_DRI_CTRL[7], Q3_LANE3_DRI_CTRL[6], 
        Q3_LANE3_DRI_CTRL[5], Q3_LANE3_DRI_CTRL[4], 
        Q3_LANE3_DRI_CTRL[3], Q3_LANE3_DRI_CTRL[2], 
        Q3_LANE3_DRI_CTRL[1], Q3_LANE3_DRI_CTRL[0]}), 
        .Q3_LANE3_DRI_RDATA({Q3_LANE3_DRI_RDATA[32], 
        Q3_LANE3_DRI_RDATA[31], Q3_LANE3_DRI_RDATA[30], 
        Q3_LANE3_DRI_RDATA[29], Q3_LANE3_DRI_RDATA[28], 
        Q3_LANE3_DRI_RDATA[27], Q3_LANE3_DRI_RDATA[26], 
        Q3_LANE3_DRI_RDATA[25], Q3_LANE3_DRI_RDATA[24], 
        Q3_LANE3_DRI_RDATA[23], Q3_LANE3_DRI_RDATA[22], 
        Q3_LANE3_DRI_RDATA[21], Q3_LANE3_DRI_RDATA[20], 
        Q3_LANE3_DRI_RDATA[19], Q3_LANE3_DRI_RDATA[18], 
        Q3_LANE3_DRI_RDATA[17], Q3_LANE3_DRI_RDATA[16], 
        Q3_LANE3_DRI_RDATA[15], Q3_LANE3_DRI_RDATA[14], 
        Q3_LANE3_DRI_RDATA[13], Q3_LANE3_DRI_RDATA[12], 
        Q3_LANE3_DRI_RDATA[11], Q3_LANE3_DRI_RDATA[10], 
        Q3_LANE3_DRI_RDATA[9], Q3_LANE3_DRI_RDATA[8], 
        Q3_LANE3_DRI_RDATA[7], Q3_LANE3_DRI_RDATA[6], 
        Q3_LANE3_DRI_RDATA[5], Q3_LANE3_DRI_RDATA[4], 
        Q3_LANE3_DRI_RDATA[3], Q3_LANE3_DRI_RDATA[2], 
        Q3_LANE3_DRI_RDATA[1], Q3_LANE3_DRI_RDATA[0]}), 
        .Q3_LANE3_DRI_INTERRUPT(Q3_LANE3_DRI_INTERRUPT), 
        .Q5_LANE0_DRI_CTRL({Q5_LANE0_DRI_CTRL[10], 
        Q5_LANE0_DRI_CTRL[9], Q5_LANE0_DRI_CTRL[8], 
        Q5_LANE0_DRI_CTRL[7], Q5_LANE0_DRI_CTRL[6], 
        Q5_LANE0_DRI_CTRL[5], Q5_LANE0_DRI_CTRL[4], 
        Q5_LANE0_DRI_CTRL[3], Q5_LANE0_DRI_CTRL[2], 
        Q5_LANE0_DRI_CTRL[1], Q5_LANE0_DRI_CTRL[0]}), 
        .Q5_LANE0_DRI_RDATA({Q5_LANE0_DRI_RDATA[32], 
        Q5_LANE0_DRI_RDATA[31], Q5_LANE0_DRI_RDATA[30], 
        Q5_LANE0_DRI_RDATA[29], Q5_LANE0_DRI_RDATA[28], 
        Q5_LANE0_DRI_RDATA[27], Q5_LANE0_DRI_RDATA[26], 
        Q5_LANE0_DRI_RDATA[25], Q5_LANE0_DRI_RDATA[24], 
        Q5_LANE0_DRI_RDATA[23], Q5_LANE0_DRI_RDATA[22], 
        Q5_LANE0_DRI_RDATA[21], Q5_LANE0_DRI_RDATA[20], 
        Q5_LANE0_DRI_RDATA[19], Q5_LANE0_DRI_RDATA[18], 
        Q5_LANE0_DRI_RDATA[17], Q5_LANE0_DRI_RDATA[16], 
        Q5_LANE0_DRI_RDATA[15], Q5_LANE0_DRI_RDATA[14], 
        Q5_LANE0_DRI_RDATA[13], Q5_LANE0_DRI_RDATA[12], 
        Q5_LANE0_DRI_RDATA[11], Q5_LANE0_DRI_RDATA[10], 
        Q5_LANE0_DRI_RDATA[9], Q5_LANE0_DRI_RDATA[8], 
        Q5_LANE0_DRI_RDATA[7], Q5_LANE0_DRI_RDATA[6], 
        Q5_LANE0_DRI_RDATA[5], Q5_LANE0_DRI_RDATA[4], 
        Q5_LANE0_DRI_RDATA[3], Q5_LANE0_DRI_RDATA[2], 
        Q5_LANE0_DRI_RDATA[1], Q5_LANE0_DRI_RDATA[0]}), 
        .Q5_LANE0_DRI_INTERRUPT(Q5_LANE0_DRI_INTERRUPT), 
        .Q5_LANE1_DRI_CTRL({Q5_LANE1_DRI_CTRL[10], 
        Q5_LANE1_DRI_CTRL[9], Q5_LANE1_DRI_CTRL[8], 
        Q5_LANE1_DRI_CTRL[7], Q5_LANE1_DRI_CTRL[6], 
        Q5_LANE1_DRI_CTRL[5], Q5_LANE1_DRI_CTRL[4], 
        Q5_LANE1_DRI_CTRL[3], Q5_LANE1_DRI_CTRL[2], 
        Q5_LANE1_DRI_CTRL[1], Q5_LANE1_DRI_CTRL[0]}), 
        .Q5_LANE1_DRI_RDATA({Q5_LANE1_DRI_RDATA[32], 
        Q5_LANE1_DRI_RDATA[31], Q5_LANE1_DRI_RDATA[30], 
        Q5_LANE1_DRI_RDATA[29], Q5_LANE1_DRI_RDATA[28], 
        Q5_LANE1_DRI_RDATA[27], Q5_LANE1_DRI_RDATA[26], 
        Q5_LANE1_DRI_RDATA[25], Q5_LANE1_DRI_RDATA[24], 
        Q5_LANE1_DRI_RDATA[23], Q5_LANE1_DRI_RDATA[22], 
        Q5_LANE1_DRI_RDATA[21], Q5_LANE1_DRI_RDATA[20], 
        Q5_LANE1_DRI_RDATA[19], Q5_LANE1_DRI_RDATA[18], 
        Q5_LANE1_DRI_RDATA[17], Q5_LANE1_DRI_RDATA[16], 
        Q5_LANE1_DRI_RDATA[15], Q5_LANE1_DRI_RDATA[14], 
        Q5_LANE1_DRI_RDATA[13], Q5_LANE1_DRI_RDATA[12], 
        Q5_LANE1_DRI_RDATA[11], Q5_LANE1_DRI_RDATA[10], 
        Q5_LANE1_DRI_RDATA[9], Q5_LANE1_DRI_RDATA[8], 
        Q5_LANE1_DRI_RDATA[7], Q5_LANE1_DRI_RDATA[6], 
        Q5_LANE1_DRI_RDATA[5], Q5_LANE1_DRI_RDATA[4], 
        Q5_LANE1_DRI_RDATA[3], Q5_LANE1_DRI_RDATA[2], 
        Q5_LANE1_DRI_RDATA[1], Q5_LANE1_DRI_RDATA[0]}), 
        .Q5_LANE1_DRI_INTERRUPT(Q5_LANE1_DRI_INTERRUPT), 
        .Q5_LANE2_DRI_CTRL({Q5_LANE2_DRI_CTRL[10], 
        Q5_LANE2_DRI_CTRL[9], Q5_LANE2_DRI_CTRL[8], 
        Q5_LANE2_DRI_CTRL[7], Q5_LANE2_DRI_CTRL[6], 
        Q5_LANE2_DRI_CTRL[5], Q5_LANE2_DRI_CTRL[4], 
        Q5_LANE2_DRI_CTRL[3], Q5_LANE2_DRI_CTRL[2], 
        Q5_LANE2_DRI_CTRL[1], Q5_LANE2_DRI_CTRL[0]}), 
        .Q5_LANE2_DRI_RDATA({Q5_LANE2_DRI_RDATA[32], 
        Q5_LANE2_DRI_RDATA[31], Q5_LANE2_DRI_RDATA[30], 
        Q5_LANE2_DRI_RDATA[29], Q5_LANE2_DRI_RDATA[28], 
        Q5_LANE2_DRI_RDATA[27], Q5_LANE2_DRI_RDATA[26], 
        Q5_LANE2_DRI_RDATA[25], Q5_LANE2_DRI_RDATA[24], 
        Q5_LANE2_DRI_RDATA[23], Q5_LANE2_DRI_RDATA[22], 
        Q5_LANE2_DRI_RDATA[21], Q5_LANE2_DRI_RDATA[20], 
        Q5_LANE2_DRI_RDATA[19], Q5_LANE2_DRI_RDATA[18], 
        Q5_LANE2_DRI_RDATA[17], Q5_LANE2_DRI_RDATA[16], 
        Q5_LANE2_DRI_RDATA[15], Q5_LANE2_DRI_RDATA[14], 
        Q5_LANE2_DRI_RDATA[13], Q5_LANE2_DRI_RDATA[12], 
        Q5_LANE2_DRI_RDATA[11], Q5_LANE2_DRI_RDATA[10], 
        Q5_LANE2_DRI_RDATA[9], Q5_LANE2_DRI_RDATA[8], 
        Q5_LANE2_DRI_RDATA[7], Q5_LANE2_DRI_RDATA[6], 
        Q5_LANE2_DRI_RDATA[5], Q5_LANE2_DRI_RDATA[4], 
        Q5_LANE2_DRI_RDATA[3], Q5_LANE2_DRI_RDATA[2], 
        Q5_LANE2_DRI_RDATA[1], Q5_LANE2_DRI_RDATA[0]}), 
        .Q5_LANE2_DRI_INTERRUPT(Q5_LANE2_DRI_INTERRUPT), 
        .Q5_LANE3_DRI_CTRL({Q5_LANE3_DRI_CTRL[10], 
        Q5_LANE3_DRI_CTRL[9], Q5_LANE3_DRI_CTRL[8], 
        Q5_LANE3_DRI_CTRL[7], Q5_LANE3_DRI_CTRL[6], 
        Q5_LANE3_DRI_CTRL[5], Q5_LANE3_DRI_CTRL[4], 
        Q5_LANE3_DRI_CTRL[3], Q5_LANE3_DRI_CTRL[2], 
        Q5_LANE3_DRI_CTRL[1], Q5_LANE3_DRI_CTRL[0]}), 
        .Q5_LANE3_DRI_RDATA({Q5_LANE3_DRI_RDATA[32], 
        Q5_LANE3_DRI_RDATA[31], Q5_LANE3_DRI_RDATA[30], 
        Q5_LANE3_DRI_RDATA[29], Q5_LANE3_DRI_RDATA[28], 
        Q5_LANE3_DRI_RDATA[27], Q5_LANE3_DRI_RDATA[26], 
        Q5_LANE3_DRI_RDATA[25], Q5_LANE3_DRI_RDATA[24], 
        Q5_LANE3_DRI_RDATA[23], Q5_LANE3_DRI_RDATA[22], 
        Q5_LANE3_DRI_RDATA[21], Q5_LANE3_DRI_RDATA[20], 
        Q5_LANE3_DRI_RDATA[19], Q5_LANE3_DRI_RDATA[18], 
        Q5_LANE3_DRI_RDATA[17], Q5_LANE3_DRI_RDATA[16], 
        Q5_LANE3_DRI_RDATA[15], Q5_LANE3_DRI_RDATA[14], 
        Q5_LANE3_DRI_RDATA[13], Q5_LANE3_DRI_RDATA[12], 
        Q5_LANE3_DRI_RDATA[11], Q5_LANE3_DRI_RDATA[10], 
        Q5_LANE3_DRI_RDATA[9], Q5_LANE3_DRI_RDATA[8], 
        Q5_LANE3_DRI_RDATA[7], Q5_LANE3_DRI_RDATA[6], 
        Q5_LANE3_DRI_RDATA[5], Q5_LANE3_DRI_RDATA[4], 
        Q5_LANE3_DRI_RDATA[3], Q5_LANE3_DRI_RDATA[2], 
        Q5_LANE3_DRI_RDATA[1], Q5_LANE3_DRI_RDATA[0]}), 
        .Q5_LANE3_DRI_INTERRUPT(Q5_LANE3_DRI_INTERRUPT), 
        .PCIE0_DRI_CTRL({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, 
        nc9, nc10}), .PCIE0_DRI_RDATA({gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net}), .PCIE0_DRI_INTERRUPT(gnd_net), 
        .PCIE1_DRI_CTRL({nc11, nc12, nc13, nc14, nc15, nc16, nc17, 
        nc18, nc19, nc20, nc21}), .PCIE1_DRI_RDATA({gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net}), .PCIE1_DRI_INTERRUPT(gnd_net), 
        .Q4_TXPLL_SSC_DRI_CTRL({Q4_TXPLL_SSC_DRI_CTRL[10], 
        Q4_TXPLL_SSC_DRI_CTRL[9], Q4_TXPLL_SSC_DRI_CTRL[8], 
        Q4_TXPLL_SSC_DRI_CTRL[7], Q4_TXPLL_SSC_DRI_CTRL[6], 
        Q4_TXPLL_SSC_DRI_CTRL[5], Q4_TXPLL_SSC_DRI_CTRL[4], 
        Q4_TXPLL_SSC_DRI_CTRL[3], Q4_TXPLL_SSC_DRI_CTRL[2], 
        Q4_TXPLL_SSC_DRI_CTRL[1], Q4_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q4_TXPLL_SSC_DRI_RDATA({Q4_TXPLL_SSC_DRI_RDATA[32], 
        Q4_TXPLL_SSC_DRI_RDATA[31], Q4_TXPLL_SSC_DRI_RDATA[30], 
        Q4_TXPLL_SSC_DRI_RDATA[29], Q4_TXPLL_SSC_DRI_RDATA[28], 
        Q4_TXPLL_SSC_DRI_RDATA[27], Q4_TXPLL_SSC_DRI_RDATA[26], 
        Q4_TXPLL_SSC_DRI_RDATA[25], Q4_TXPLL_SSC_DRI_RDATA[24], 
        Q4_TXPLL_SSC_DRI_RDATA[23], Q4_TXPLL_SSC_DRI_RDATA[22], 
        Q4_TXPLL_SSC_DRI_RDATA[21], Q4_TXPLL_SSC_DRI_RDATA[20], 
        Q4_TXPLL_SSC_DRI_RDATA[19], Q4_TXPLL_SSC_DRI_RDATA[18], 
        Q4_TXPLL_SSC_DRI_RDATA[17], Q4_TXPLL_SSC_DRI_RDATA[16], 
        Q4_TXPLL_SSC_DRI_RDATA[15], Q4_TXPLL_SSC_DRI_RDATA[14], 
        Q4_TXPLL_SSC_DRI_RDATA[13], Q4_TXPLL_SSC_DRI_RDATA[12], 
        Q4_TXPLL_SSC_DRI_RDATA[11], Q4_TXPLL_SSC_DRI_RDATA[10], 
        Q4_TXPLL_SSC_DRI_RDATA[9], Q4_TXPLL_SSC_DRI_RDATA[8], 
        Q4_TXPLL_SSC_DRI_RDATA[7], Q4_TXPLL_SSC_DRI_RDATA[6], 
        Q4_TXPLL_SSC_DRI_RDATA[5], Q4_TXPLL_SSC_DRI_RDATA[4], 
        Q4_TXPLL_SSC_DRI_RDATA[3], Q4_TXPLL_SSC_DRI_RDATA[2], 
        Q4_TXPLL_SSC_DRI_RDATA[1], Q4_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q4_TXPLL_SSC_DRI_INTERRUPT(Q4_TXPLL_SSC_DRI_INTERRUPT), 
        .Q2_TXPLL_SSC_DRI_CTRL({Q2_TXPLL_SSC_DRI_CTRL[10], 
        Q2_TXPLL_SSC_DRI_CTRL[9], Q2_TXPLL_SSC_DRI_CTRL[8], 
        Q2_TXPLL_SSC_DRI_CTRL[7], Q2_TXPLL_SSC_DRI_CTRL[6], 
        Q2_TXPLL_SSC_DRI_CTRL[5], Q2_TXPLL_SSC_DRI_CTRL[4], 
        Q2_TXPLL_SSC_DRI_CTRL[3], Q2_TXPLL_SSC_DRI_CTRL[2], 
        Q2_TXPLL_SSC_DRI_CTRL[1], Q2_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q2_TXPLL_SSC_DRI_RDATA({Q2_TXPLL_SSC_DRI_RDATA[32], 
        Q2_TXPLL_SSC_DRI_RDATA[31], Q2_TXPLL_SSC_DRI_RDATA[30], 
        Q2_TXPLL_SSC_DRI_RDATA[29], Q2_TXPLL_SSC_DRI_RDATA[28], 
        Q2_TXPLL_SSC_DRI_RDATA[27], Q2_TXPLL_SSC_DRI_RDATA[26], 
        Q2_TXPLL_SSC_DRI_RDATA[25], Q2_TXPLL_SSC_DRI_RDATA[24], 
        Q2_TXPLL_SSC_DRI_RDATA[23], Q2_TXPLL_SSC_DRI_RDATA[22], 
        Q2_TXPLL_SSC_DRI_RDATA[21], Q2_TXPLL_SSC_DRI_RDATA[20], 
        Q2_TXPLL_SSC_DRI_RDATA[19], Q2_TXPLL_SSC_DRI_RDATA[18], 
        Q2_TXPLL_SSC_DRI_RDATA[17], Q2_TXPLL_SSC_DRI_RDATA[16], 
        Q2_TXPLL_SSC_DRI_RDATA[15], Q2_TXPLL_SSC_DRI_RDATA[14], 
        Q2_TXPLL_SSC_DRI_RDATA[13], Q2_TXPLL_SSC_DRI_RDATA[12], 
        Q2_TXPLL_SSC_DRI_RDATA[11], Q2_TXPLL_SSC_DRI_RDATA[10], 
        Q2_TXPLL_SSC_DRI_RDATA[9], Q2_TXPLL_SSC_DRI_RDATA[8], 
        Q2_TXPLL_SSC_DRI_RDATA[7], Q2_TXPLL_SSC_DRI_RDATA[6], 
        Q2_TXPLL_SSC_DRI_RDATA[5], Q2_TXPLL_SSC_DRI_RDATA[4], 
        Q2_TXPLL_SSC_DRI_RDATA[3], Q2_TXPLL_SSC_DRI_RDATA[2], 
        Q2_TXPLL_SSC_DRI_RDATA[1], Q2_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q2_TXPLL_SSC_DRI_INTERRUPT(Q2_TXPLL_SSC_DRI_INTERRUPT), 
        .Q0_TXPLL_SSC_DRI_CTRL({Q0_TXPLL_SSC_DRI_CTRL[10], 
        Q0_TXPLL_SSC_DRI_CTRL[9], Q0_TXPLL_SSC_DRI_CTRL[8], 
        Q0_TXPLL_SSC_DRI_CTRL[7], Q0_TXPLL_SSC_DRI_CTRL[6], 
        Q0_TXPLL_SSC_DRI_CTRL[5], Q0_TXPLL_SSC_DRI_CTRL[4], 
        Q0_TXPLL_SSC_DRI_CTRL[3], Q0_TXPLL_SSC_DRI_CTRL[2], 
        Q0_TXPLL_SSC_DRI_CTRL[1], Q0_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q0_TXPLL_SSC_DRI_RDATA({Q0_TXPLL_SSC_DRI_RDATA[32], 
        Q0_TXPLL_SSC_DRI_RDATA[31], Q0_TXPLL_SSC_DRI_RDATA[30], 
        Q0_TXPLL_SSC_DRI_RDATA[29], Q0_TXPLL_SSC_DRI_RDATA[28], 
        Q0_TXPLL_SSC_DRI_RDATA[27], Q0_TXPLL_SSC_DRI_RDATA[26], 
        Q0_TXPLL_SSC_DRI_RDATA[25], Q0_TXPLL_SSC_DRI_RDATA[24], 
        Q0_TXPLL_SSC_DRI_RDATA[23], Q0_TXPLL_SSC_DRI_RDATA[22], 
        Q0_TXPLL_SSC_DRI_RDATA[21], Q0_TXPLL_SSC_DRI_RDATA[20], 
        Q0_TXPLL_SSC_DRI_RDATA[19], Q0_TXPLL_SSC_DRI_RDATA[18], 
        Q0_TXPLL_SSC_DRI_RDATA[17], Q0_TXPLL_SSC_DRI_RDATA[16], 
        Q0_TXPLL_SSC_DRI_RDATA[15], Q0_TXPLL_SSC_DRI_RDATA[14], 
        Q0_TXPLL_SSC_DRI_RDATA[13], Q0_TXPLL_SSC_DRI_RDATA[12], 
        Q0_TXPLL_SSC_DRI_RDATA[11], Q0_TXPLL_SSC_DRI_RDATA[10], 
        Q0_TXPLL_SSC_DRI_RDATA[9], Q0_TXPLL_SSC_DRI_RDATA[8], 
        Q0_TXPLL_SSC_DRI_RDATA[7], Q0_TXPLL_SSC_DRI_RDATA[6], 
        Q0_TXPLL_SSC_DRI_RDATA[5], Q0_TXPLL_SSC_DRI_RDATA[4], 
        Q0_TXPLL_SSC_DRI_RDATA[3], Q0_TXPLL_SSC_DRI_RDATA[2], 
        Q0_TXPLL_SSC_DRI_RDATA[1], Q0_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q0_TXPLL_SSC_DRI_INTERRUPT(Q0_TXPLL_SSC_DRI_INTERRUPT), 
        .Q1_TXPLL_SSC_DRI_CTRL({Q1_TXPLL_SSC_DRI_CTRL[10], 
        Q1_TXPLL_SSC_DRI_CTRL[9], Q1_TXPLL_SSC_DRI_CTRL[8], 
        Q1_TXPLL_SSC_DRI_CTRL[7], Q1_TXPLL_SSC_DRI_CTRL[6], 
        Q1_TXPLL_SSC_DRI_CTRL[5], Q1_TXPLL_SSC_DRI_CTRL[4], 
        Q1_TXPLL_SSC_DRI_CTRL[3], Q1_TXPLL_SSC_DRI_CTRL[2], 
        Q1_TXPLL_SSC_DRI_CTRL[1], Q1_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q1_TXPLL_SSC_DRI_RDATA({Q1_TXPLL_SSC_DRI_RDATA[32], 
        Q1_TXPLL_SSC_DRI_RDATA[31], Q1_TXPLL_SSC_DRI_RDATA[30], 
        Q1_TXPLL_SSC_DRI_RDATA[29], Q1_TXPLL_SSC_DRI_RDATA[28], 
        Q1_TXPLL_SSC_DRI_RDATA[27], Q1_TXPLL_SSC_DRI_RDATA[26], 
        Q1_TXPLL_SSC_DRI_RDATA[25], Q1_TXPLL_SSC_DRI_RDATA[24], 
        Q1_TXPLL_SSC_DRI_RDATA[23], Q1_TXPLL_SSC_DRI_RDATA[22], 
        Q1_TXPLL_SSC_DRI_RDATA[21], Q1_TXPLL_SSC_DRI_RDATA[20], 
        Q1_TXPLL_SSC_DRI_RDATA[19], Q1_TXPLL_SSC_DRI_RDATA[18], 
        Q1_TXPLL_SSC_DRI_RDATA[17], Q1_TXPLL_SSC_DRI_RDATA[16], 
        Q1_TXPLL_SSC_DRI_RDATA[15], Q1_TXPLL_SSC_DRI_RDATA[14], 
        Q1_TXPLL_SSC_DRI_RDATA[13], Q1_TXPLL_SSC_DRI_RDATA[12], 
        Q1_TXPLL_SSC_DRI_RDATA[11], Q1_TXPLL_SSC_DRI_RDATA[10], 
        Q1_TXPLL_SSC_DRI_RDATA[9], Q1_TXPLL_SSC_DRI_RDATA[8], 
        Q1_TXPLL_SSC_DRI_RDATA[7], Q1_TXPLL_SSC_DRI_RDATA[6], 
        Q1_TXPLL_SSC_DRI_RDATA[5], Q1_TXPLL_SSC_DRI_RDATA[4], 
        Q1_TXPLL_SSC_DRI_RDATA[3], Q1_TXPLL_SSC_DRI_RDATA[2], 
        Q1_TXPLL_SSC_DRI_RDATA[1], Q1_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q1_TXPLL_SSC_DRI_INTERRUPT(Q1_TXPLL_SSC_DRI_INTERRUPT), 
        .Q3_TXPLL_SSC_DRI_CTRL({Q3_TXPLL_SSC_DRI_CTRL[10], 
        Q3_TXPLL_SSC_DRI_CTRL[9], Q3_TXPLL_SSC_DRI_CTRL[8], 
        Q3_TXPLL_SSC_DRI_CTRL[7], Q3_TXPLL_SSC_DRI_CTRL[6], 
        Q3_TXPLL_SSC_DRI_CTRL[5], Q3_TXPLL_SSC_DRI_CTRL[4], 
        Q3_TXPLL_SSC_DRI_CTRL[3], Q3_TXPLL_SSC_DRI_CTRL[2], 
        Q3_TXPLL_SSC_DRI_CTRL[1], Q3_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q3_TXPLL_SSC_DRI_RDATA({Q3_TXPLL_SSC_DRI_RDATA[32], 
        Q3_TXPLL_SSC_DRI_RDATA[31], Q3_TXPLL_SSC_DRI_RDATA[30], 
        Q3_TXPLL_SSC_DRI_RDATA[29], Q3_TXPLL_SSC_DRI_RDATA[28], 
        Q3_TXPLL_SSC_DRI_RDATA[27], Q3_TXPLL_SSC_DRI_RDATA[26], 
        Q3_TXPLL_SSC_DRI_RDATA[25], Q3_TXPLL_SSC_DRI_RDATA[24], 
        Q3_TXPLL_SSC_DRI_RDATA[23], Q3_TXPLL_SSC_DRI_RDATA[22], 
        Q3_TXPLL_SSC_DRI_RDATA[21], Q3_TXPLL_SSC_DRI_RDATA[20], 
        Q3_TXPLL_SSC_DRI_RDATA[19], Q3_TXPLL_SSC_DRI_RDATA[18], 
        Q3_TXPLL_SSC_DRI_RDATA[17], Q3_TXPLL_SSC_DRI_RDATA[16], 
        Q3_TXPLL_SSC_DRI_RDATA[15], Q3_TXPLL_SSC_DRI_RDATA[14], 
        Q3_TXPLL_SSC_DRI_RDATA[13], Q3_TXPLL_SSC_DRI_RDATA[12], 
        Q3_TXPLL_SSC_DRI_RDATA[11], Q3_TXPLL_SSC_DRI_RDATA[10], 
        Q3_TXPLL_SSC_DRI_RDATA[9], Q3_TXPLL_SSC_DRI_RDATA[8], 
        Q3_TXPLL_SSC_DRI_RDATA[7], Q3_TXPLL_SSC_DRI_RDATA[6], 
        Q3_TXPLL_SSC_DRI_RDATA[5], Q3_TXPLL_SSC_DRI_RDATA[4], 
        Q3_TXPLL_SSC_DRI_RDATA[3], Q3_TXPLL_SSC_DRI_RDATA[2], 
        Q3_TXPLL_SSC_DRI_RDATA[1], Q3_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q3_TXPLL_SSC_DRI_INTERRUPT(Q3_TXPLL_SSC_DRI_INTERRUPT), 
        .Q5_TXPLL_SSC_DRI_CTRL({Q5_TXPLL_SSC_DRI_CTRL[10], 
        Q5_TXPLL_SSC_DRI_CTRL[9], Q5_TXPLL_SSC_DRI_CTRL[8], 
        Q5_TXPLL_SSC_DRI_CTRL[7], Q5_TXPLL_SSC_DRI_CTRL[6], 
        Q5_TXPLL_SSC_DRI_CTRL[5], Q5_TXPLL_SSC_DRI_CTRL[4], 
        Q5_TXPLL_SSC_DRI_CTRL[3], Q5_TXPLL_SSC_DRI_CTRL[2], 
        Q5_TXPLL_SSC_DRI_CTRL[1], Q5_TXPLL_SSC_DRI_CTRL[0]}), 
        .Q5_TXPLL_SSC_DRI_RDATA({Q5_TXPLL_SSC_DRI_RDATA[32], 
        Q5_TXPLL_SSC_DRI_RDATA[31], Q5_TXPLL_SSC_DRI_RDATA[30], 
        Q5_TXPLL_SSC_DRI_RDATA[29], Q5_TXPLL_SSC_DRI_RDATA[28], 
        Q5_TXPLL_SSC_DRI_RDATA[27], Q5_TXPLL_SSC_DRI_RDATA[26], 
        Q5_TXPLL_SSC_DRI_RDATA[25], Q5_TXPLL_SSC_DRI_RDATA[24], 
        Q5_TXPLL_SSC_DRI_RDATA[23], Q5_TXPLL_SSC_DRI_RDATA[22], 
        Q5_TXPLL_SSC_DRI_RDATA[21], Q5_TXPLL_SSC_DRI_RDATA[20], 
        Q5_TXPLL_SSC_DRI_RDATA[19], Q5_TXPLL_SSC_DRI_RDATA[18], 
        Q5_TXPLL_SSC_DRI_RDATA[17], Q5_TXPLL_SSC_DRI_RDATA[16], 
        Q5_TXPLL_SSC_DRI_RDATA[15], Q5_TXPLL_SSC_DRI_RDATA[14], 
        Q5_TXPLL_SSC_DRI_RDATA[13], Q5_TXPLL_SSC_DRI_RDATA[12], 
        Q5_TXPLL_SSC_DRI_RDATA[11], Q5_TXPLL_SSC_DRI_RDATA[10], 
        Q5_TXPLL_SSC_DRI_RDATA[9], Q5_TXPLL_SSC_DRI_RDATA[8], 
        Q5_TXPLL_SSC_DRI_RDATA[7], Q5_TXPLL_SSC_DRI_RDATA[6], 
        Q5_TXPLL_SSC_DRI_RDATA[5], Q5_TXPLL_SSC_DRI_RDATA[4], 
        Q5_TXPLL_SSC_DRI_RDATA[3], Q5_TXPLL_SSC_DRI_RDATA[2], 
        Q5_TXPLL_SSC_DRI_RDATA[1], Q5_TXPLL_SSC_DRI_RDATA[0]}), 
        .Q5_TXPLL_SSC_DRI_INTERRUPT(Q5_TXPLL_SSC_DRI_INTERRUPT), 
        .Q4_TXPLL_DRI_CTRL({Q4_TXPLL_DRI_CTRL[10], 
        Q4_TXPLL_DRI_CTRL[9], Q4_TXPLL_DRI_CTRL[8], 
        Q4_TXPLL_DRI_CTRL[7], Q4_TXPLL_DRI_CTRL[6], 
        Q4_TXPLL_DRI_CTRL[5], Q4_TXPLL_DRI_CTRL[4], 
        Q4_TXPLL_DRI_CTRL[3], Q4_TXPLL_DRI_CTRL[2], 
        Q4_TXPLL_DRI_CTRL[1], Q4_TXPLL_DRI_CTRL[0]}), 
        .Q4_TXPLL_DRI_RDATA({Q4_TXPLL_DRI_RDATA[32], 
        Q4_TXPLL_DRI_RDATA[31], Q4_TXPLL_DRI_RDATA[30], 
        Q4_TXPLL_DRI_RDATA[29], Q4_TXPLL_DRI_RDATA[28], 
        Q4_TXPLL_DRI_RDATA[27], Q4_TXPLL_DRI_RDATA[26], 
        Q4_TXPLL_DRI_RDATA[25], Q4_TXPLL_DRI_RDATA[24], 
        Q4_TXPLL_DRI_RDATA[23], Q4_TXPLL_DRI_RDATA[22], 
        Q4_TXPLL_DRI_RDATA[21], Q4_TXPLL_DRI_RDATA[20], 
        Q4_TXPLL_DRI_RDATA[19], Q4_TXPLL_DRI_RDATA[18], 
        Q4_TXPLL_DRI_RDATA[17], Q4_TXPLL_DRI_RDATA[16], 
        Q4_TXPLL_DRI_RDATA[15], Q4_TXPLL_DRI_RDATA[14], 
        Q4_TXPLL_DRI_RDATA[13], Q4_TXPLL_DRI_RDATA[12], 
        Q4_TXPLL_DRI_RDATA[11], Q4_TXPLL_DRI_RDATA[10], 
        Q4_TXPLL_DRI_RDATA[9], Q4_TXPLL_DRI_RDATA[8], 
        Q4_TXPLL_DRI_RDATA[7], Q4_TXPLL_DRI_RDATA[6], 
        Q4_TXPLL_DRI_RDATA[5], Q4_TXPLL_DRI_RDATA[4], 
        Q4_TXPLL_DRI_RDATA[3], Q4_TXPLL_DRI_RDATA[2], 
        Q4_TXPLL_DRI_RDATA[1], Q4_TXPLL_DRI_RDATA[0]}), 
        .Q4_TXPLL_DRI_INTERRUPT(Q4_TXPLL_DRI_INTERRUPT), 
        .Q2_TXPLL0_DRI_CTRL({Q2_TXPLL0_DRI_CTRL[10], 
        Q2_TXPLL0_DRI_CTRL[9], Q2_TXPLL0_DRI_CTRL[8], 
        Q2_TXPLL0_DRI_CTRL[7], Q2_TXPLL0_DRI_CTRL[6], 
        Q2_TXPLL0_DRI_CTRL[5], Q2_TXPLL0_DRI_CTRL[4], 
        Q2_TXPLL0_DRI_CTRL[3], Q2_TXPLL0_DRI_CTRL[2], 
        Q2_TXPLL0_DRI_CTRL[1], Q2_TXPLL0_DRI_CTRL[0]}), 
        .Q2_TXPLL0_DRI_RDATA({Q2_TXPLL0_DRI_RDATA[32], 
        Q2_TXPLL0_DRI_RDATA[31], Q2_TXPLL0_DRI_RDATA[30], 
        Q2_TXPLL0_DRI_RDATA[29], Q2_TXPLL0_DRI_RDATA[28], 
        Q2_TXPLL0_DRI_RDATA[27], Q2_TXPLL0_DRI_RDATA[26], 
        Q2_TXPLL0_DRI_RDATA[25], Q2_TXPLL0_DRI_RDATA[24], 
        Q2_TXPLL0_DRI_RDATA[23], Q2_TXPLL0_DRI_RDATA[22], 
        Q2_TXPLL0_DRI_RDATA[21], Q2_TXPLL0_DRI_RDATA[20], 
        Q2_TXPLL0_DRI_RDATA[19], Q2_TXPLL0_DRI_RDATA[18], 
        Q2_TXPLL0_DRI_RDATA[17], Q2_TXPLL0_DRI_RDATA[16], 
        Q2_TXPLL0_DRI_RDATA[15], Q2_TXPLL0_DRI_RDATA[14], 
        Q2_TXPLL0_DRI_RDATA[13], Q2_TXPLL0_DRI_RDATA[12], 
        Q2_TXPLL0_DRI_RDATA[11], Q2_TXPLL0_DRI_RDATA[10], 
        Q2_TXPLL0_DRI_RDATA[9], Q2_TXPLL0_DRI_RDATA[8], 
        Q2_TXPLL0_DRI_RDATA[7], Q2_TXPLL0_DRI_RDATA[6], 
        Q2_TXPLL0_DRI_RDATA[5], Q2_TXPLL0_DRI_RDATA[4], 
        Q2_TXPLL0_DRI_RDATA[3], Q2_TXPLL0_DRI_RDATA[2], 
        Q2_TXPLL0_DRI_RDATA[1], Q2_TXPLL0_DRI_RDATA[0]}), 
        .Q2_TXPLL0_DRI_INTERRUPT(Q2_TXPLL0_DRI_INTERRUPT), 
        .Q2_TXPLL1_DRI_CTRL({Q2_TXPLL1_DRI_CTRL[10], 
        Q2_TXPLL1_DRI_CTRL[9], Q2_TXPLL1_DRI_CTRL[8], 
        Q2_TXPLL1_DRI_CTRL[7], Q2_TXPLL1_DRI_CTRL[6], 
        Q2_TXPLL1_DRI_CTRL[5], Q2_TXPLL1_DRI_CTRL[4], 
        Q2_TXPLL1_DRI_CTRL[3], Q2_TXPLL1_DRI_CTRL[2], 
        Q2_TXPLL1_DRI_CTRL[1], Q2_TXPLL1_DRI_CTRL[0]}), 
        .Q2_TXPLL1_DRI_RDATA({Q2_TXPLL1_DRI_RDATA[32], 
        Q2_TXPLL1_DRI_RDATA[31], Q2_TXPLL1_DRI_RDATA[30], 
        Q2_TXPLL1_DRI_RDATA[29], Q2_TXPLL1_DRI_RDATA[28], 
        Q2_TXPLL1_DRI_RDATA[27], Q2_TXPLL1_DRI_RDATA[26], 
        Q2_TXPLL1_DRI_RDATA[25], Q2_TXPLL1_DRI_RDATA[24], 
        Q2_TXPLL1_DRI_RDATA[23], Q2_TXPLL1_DRI_RDATA[22], 
        Q2_TXPLL1_DRI_RDATA[21], Q2_TXPLL1_DRI_RDATA[20], 
        Q2_TXPLL1_DRI_RDATA[19], Q2_TXPLL1_DRI_RDATA[18], 
        Q2_TXPLL1_DRI_RDATA[17], Q2_TXPLL1_DRI_RDATA[16], 
        Q2_TXPLL1_DRI_RDATA[15], Q2_TXPLL1_DRI_RDATA[14], 
        Q2_TXPLL1_DRI_RDATA[13], Q2_TXPLL1_DRI_RDATA[12], 
        Q2_TXPLL1_DRI_RDATA[11], Q2_TXPLL1_DRI_RDATA[10], 
        Q2_TXPLL1_DRI_RDATA[9], Q2_TXPLL1_DRI_RDATA[8], 
        Q2_TXPLL1_DRI_RDATA[7], Q2_TXPLL1_DRI_RDATA[6], 
        Q2_TXPLL1_DRI_RDATA[5], Q2_TXPLL1_DRI_RDATA[4], 
        Q2_TXPLL1_DRI_RDATA[3], Q2_TXPLL1_DRI_RDATA[2], 
        Q2_TXPLL1_DRI_RDATA[1], Q2_TXPLL1_DRI_RDATA[0]}), 
        .Q2_TXPLL1_DRI_INTERRUPT(Q2_TXPLL1_DRI_INTERRUPT), 
        .Q0_TXPLL0_DRI_CTRL({Q0_TXPLL0_DRI_CTRL[10], 
        Q0_TXPLL0_DRI_CTRL[9], Q0_TXPLL0_DRI_CTRL[8], 
        Q0_TXPLL0_DRI_CTRL[7], Q0_TXPLL0_DRI_CTRL[6], 
        Q0_TXPLL0_DRI_CTRL[5], Q0_TXPLL0_DRI_CTRL[4], 
        Q0_TXPLL0_DRI_CTRL[3], Q0_TXPLL0_DRI_CTRL[2], 
        Q0_TXPLL0_DRI_CTRL[1], Q0_TXPLL0_DRI_CTRL[0]}), 
        .Q0_TXPLL0_DRI_RDATA({Q0_TXPLL0_DRI_RDATA[32], 
        Q0_TXPLL0_DRI_RDATA[31], Q0_TXPLL0_DRI_RDATA[30], 
        Q0_TXPLL0_DRI_RDATA[29], Q0_TXPLL0_DRI_RDATA[28], 
        Q0_TXPLL0_DRI_RDATA[27], Q0_TXPLL0_DRI_RDATA[26], 
        Q0_TXPLL0_DRI_RDATA[25], Q0_TXPLL0_DRI_RDATA[24], 
        Q0_TXPLL0_DRI_RDATA[23], Q0_TXPLL0_DRI_RDATA[22], 
        Q0_TXPLL0_DRI_RDATA[21], Q0_TXPLL0_DRI_RDATA[20], 
        Q0_TXPLL0_DRI_RDATA[19], Q0_TXPLL0_DRI_RDATA[18], 
        Q0_TXPLL0_DRI_RDATA[17], Q0_TXPLL0_DRI_RDATA[16], 
        Q0_TXPLL0_DRI_RDATA[15], Q0_TXPLL0_DRI_RDATA[14], 
        Q0_TXPLL0_DRI_RDATA[13], Q0_TXPLL0_DRI_RDATA[12], 
        Q0_TXPLL0_DRI_RDATA[11], Q0_TXPLL0_DRI_RDATA[10], 
        Q0_TXPLL0_DRI_RDATA[9], Q0_TXPLL0_DRI_RDATA[8], 
        Q0_TXPLL0_DRI_RDATA[7], Q0_TXPLL0_DRI_RDATA[6], 
        Q0_TXPLL0_DRI_RDATA[5], Q0_TXPLL0_DRI_RDATA[4], 
        Q0_TXPLL0_DRI_RDATA[3], Q0_TXPLL0_DRI_RDATA[2], 
        Q0_TXPLL0_DRI_RDATA[1], Q0_TXPLL0_DRI_RDATA[0]}), 
        .Q0_TXPLL0_DRI_INTERRUPT(Q0_TXPLL0_DRI_INTERRUPT), 
        .Q0_TXPLL1_DRI_CTRL({Q0_TXPLL1_DRI_CTRL[10], 
        Q0_TXPLL1_DRI_CTRL[9], Q0_TXPLL1_DRI_CTRL[8], 
        Q0_TXPLL1_DRI_CTRL[7], Q0_TXPLL1_DRI_CTRL[6], 
        Q0_TXPLL1_DRI_CTRL[5], Q0_TXPLL1_DRI_CTRL[4], 
        Q0_TXPLL1_DRI_CTRL[3], Q0_TXPLL1_DRI_CTRL[2], 
        Q0_TXPLL1_DRI_CTRL[1], Q0_TXPLL1_DRI_CTRL[0]}), 
        .Q0_TXPLL1_DRI_RDATA({Q0_TXPLL1_DRI_RDATA[32], 
        Q0_TXPLL1_DRI_RDATA[31], Q0_TXPLL1_DRI_RDATA[30], 
        Q0_TXPLL1_DRI_RDATA[29], Q0_TXPLL1_DRI_RDATA[28], 
        Q0_TXPLL1_DRI_RDATA[27], Q0_TXPLL1_DRI_RDATA[26], 
        Q0_TXPLL1_DRI_RDATA[25], Q0_TXPLL1_DRI_RDATA[24], 
        Q0_TXPLL1_DRI_RDATA[23], Q0_TXPLL1_DRI_RDATA[22], 
        Q0_TXPLL1_DRI_RDATA[21], Q0_TXPLL1_DRI_RDATA[20], 
        Q0_TXPLL1_DRI_RDATA[19], Q0_TXPLL1_DRI_RDATA[18], 
        Q0_TXPLL1_DRI_RDATA[17], Q0_TXPLL1_DRI_RDATA[16], 
        Q0_TXPLL1_DRI_RDATA[15], Q0_TXPLL1_DRI_RDATA[14], 
        Q0_TXPLL1_DRI_RDATA[13], Q0_TXPLL1_DRI_RDATA[12], 
        Q0_TXPLL1_DRI_RDATA[11], Q0_TXPLL1_DRI_RDATA[10], 
        Q0_TXPLL1_DRI_RDATA[9], Q0_TXPLL1_DRI_RDATA[8], 
        Q0_TXPLL1_DRI_RDATA[7], Q0_TXPLL1_DRI_RDATA[6], 
        Q0_TXPLL1_DRI_RDATA[5], Q0_TXPLL1_DRI_RDATA[4], 
        Q0_TXPLL1_DRI_RDATA[3], Q0_TXPLL1_DRI_RDATA[2], 
        Q0_TXPLL1_DRI_RDATA[1], Q0_TXPLL1_DRI_RDATA[0]}), 
        .Q0_TXPLL1_DRI_INTERRUPT(Q0_TXPLL1_DRI_INTERRUPT), 
        .Q1_TXPLL0_DRI_CTRL({Q1_TXPLL0_DRI_CTRL[10], 
        Q1_TXPLL0_DRI_CTRL[9], Q1_TXPLL0_DRI_CTRL[8], 
        Q1_TXPLL0_DRI_CTRL[7], Q1_TXPLL0_DRI_CTRL[6], 
        Q1_TXPLL0_DRI_CTRL[5], Q1_TXPLL0_DRI_CTRL[4], 
        Q1_TXPLL0_DRI_CTRL[3], Q1_TXPLL0_DRI_CTRL[2], 
        Q1_TXPLL0_DRI_CTRL[1], Q1_TXPLL0_DRI_CTRL[0]}), 
        .Q1_TXPLL0_DRI_RDATA({Q1_TXPLL0_DRI_RDATA[32], 
        Q1_TXPLL0_DRI_RDATA[31], Q1_TXPLL0_DRI_RDATA[30], 
        Q1_TXPLL0_DRI_RDATA[29], Q1_TXPLL0_DRI_RDATA[28], 
        Q1_TXPLL0_DRI_RDATA[27], Q1_TXPLL0_DRI_RDATA[26], 
        Q1_TXPLL0_DRI_RDATA[25], Q1_TXPLL0_DRI_RDATA[24], 
        Q1_TXPLL0_DRI_RDATA[23], Q1_TXPLL0_DRI_RDATA[22], 
        Q1_TXPLL0_DRI_RDATA[21], Q1_TXPLL0_DRI_RDATA[20], 
        Q1_TXPLL0_DRI_RDATA[19], Q1_TXPLL0_DRI_RDATA[18], 
        Q1_TXPLL0_DRI_RDATA[17], Q1_TXPLL0_DRI_RDATA[16], 
        Q1_TXPLL0_DRI_RDATA[15], Q1_TXPLL0_DRI_RDATA[14], 
        Q1_TXPLL0_DRI_RDATA[13], Q1_TXPLL0_DRI_RDATA[12], 
        Q1_TXPLL0_DRI_RDATA[11], Q1_TXPLL0_DRI_RDATA[10], 
        Q1_TXPLL0_DRI_RDATA[9], Q1_TXPLL0_DRI_RDATA[8], 
        Q1_TXPLL0_DRI_RDATA[7], Q1_TXPLL0_DRI_RDATA[6], 
        Q1_TXPLL0_DRI_RDATA[5], Q1_TXPLL0_DRI_RDATA[4], 
        Q1_TXPLL0_DRI_RDATA[3], Q1_TXPLL0_DRI_RDATA[2], 
        Q1_TXPLL0_DRI_RDATA[1], Q1_TXPLL0_DRI_RDATA[0]}), 
        .Q1_TXPLL0_DRI_INTERRUPT(Q1_TXPLL0_DRI_INTERRUPT), 
        .Q1_TXPLL1_DRI_CTRL({Q1_TXPLL1_DRI_CTRL[10], 
        Q1_TXPLL1_DRI_CTRL[9], Q1_TXPLL1_DRI_CTRL[8], 
        Q1_TXPLL1_DRI_CTRL[7], Q1_TXPLL1_DRI_CTRL[6], 
        Q1_TXPLL1_DRI_CTRL[5], Q1_TXPLL1_DRI_CTRL[4], 
        Q1_TXPLL1_DRI_CTRL[3], Q1_TXPLL1_DRI_CTRL[2], 
        Q1_TXPLL1_DRI_CTRL[1], Q1_TXPLL1_DRI_CTRL[0]}), 
        .Q1_TXPLL1_DRI_RDATA({Q1_TXPLL1_DRI_RDATA[32], 
        Q1_TXPLL1_DRI_RDATA[31], Q1_TXPLL1_DRI_RDATA[30], 
        Q1_TXPLL1_DRI_RDATA[29], Q1_TXPLL1_DRI_RDATA[28], 
        Q1_TXPLL1_DRI_RDATA[27], Q1_TXPLL1_DRI_RDATA[26], 
        Q1_TXPLL1_DRI_RDATA[25], Q1_TXPLL1_DRI_RDATA[24], 
        Q1_TXPLL1_DRI_RDATA[23], Q1_TXPLL1_DRI_RDATA[22], 
        Q1_TXPLL1_DRI_RDATA[21], Q1_TXPLL1_DRI_RDATA[20], 
        Q1_TXPLL1_DRI_RDATA[19], Q1_TXPLL1_DRI_RDATA[18], 
        Q1_TXPLL1_DRI_RDATA[17], Q1_TXPLL1_DRI_RDATA[16], 
        Q1_TXPLL1_DRI_RDATA[15], Q1_TXPLL1_DRI_RDATA[14], 
        Q1_TXPLL1_DRI_RDATA[13], Q1_TXPLL1_DRI_RDATA[12], 
        Q1_TXPLL1_DRI_RDATA[11], Q1_TXPLL1_DRI_RDATA[10], 
        Q1_TXPLL1_DRI_RDATA[9], Q1_TXPLL1_DRI_RDATA[8], 
        Q1_TXPLL1_DRI_RDATA[7], Q1_TXPLL1_DRI_RDATA[6], 
        Q1_TXPLL1_DRI_RDATA[5], Q1_TXPLL1_DRI_RDATA[4], 
        Q1_TXPLL1_DRI_RDATA[3], Q1_TXPLL1_DRI_RDATA[2], 
        Q1_TXPLL1_DRI_RDATA[1], Q1_TXPLL1_DRI_RDATA[0]}), 
        .Q1_TXPLL1_DRI_INTERRUPT(Q1_TXPLL1_DRI_INTERRUPT), 
        .Q3_TXPLL_DRI_CTRL({Q3_TXPLL_DRI_CTRL[10], 
        Q3_TXPLL_DRI_CTRL[9], Q3_TXPLL_DRI_CTRL[8], 
        Q3_TXPLL_DRI_CTRL[7], Q3_TXPLL_DRI_CTRL[6], 
        Q3_TXPLL_DRI_CTRL[5], Q3_TXPLL_DRI_CTRL[4], 
        Q3_TXPLL_DRI_CTRL[3], Q3_TXPLL_DRI_CTRL[2], 
        Q3_TXPLL_DRI_CTRL[1], Q3_TXPLL_DRI_CTRL[0]}), 
        .Q3_TXPLL_DRI_RDATA({Q3_TXPLL_DRI_RDATA[32], 
        Q3_TXPLL_DRI_RDATA[31], Q3_TXPLL_DRI_RDATA[30], 
        Q3_TXPLL_DRI_RDATA[29], Q3_TXPLL_DRI_RDATA[28], 
        Q3_TXPLL_DRI_RDATA[27], Q3_TXPLL_DRI_RDATA[26], 
        Q3_TXPLL_DRI_RDATA[25], Q3_TXPLL_DRI_RDATA[24], 
        Q3_TXPLL_DRI_RDATA[23], Q3_TXPLL_DRI_RDATA[22], 
        Q3_TXPLL_DRI_RDATA[21], Q3_TXPLL_DRI_RDATA[20], 
        Q3_TXPLL_DRI_RDATA[19], Q3_TXPLL_DRI_RDATA[18], 
        Q3_TXPLL_DRI_RDATA[17], Q3_TXPLL_DRI_RDATA[16], 
        Q3_TXPLL_DRI_RDATA[15], Q3_TXPLL_DRI_RDATA[14], 
        Q3_TXPLL_DRI_RDATA[13], Q3_TXPLL_DRI_RDATA[12], 
        Q3_TXPLL_DRI_RDATA[11], Q3_TXPLL_DRI_RDATA[10], 
        Q3_TXPLL_DRI_RDATA[9], Q3_TXPLL_DRI_RDATA[8], 
        Q3_TXPLL_DRI_RDATA[7], Q3_TXPLL_DRI_RDATA[6], 
        Q3_TXPLL_DRI_RDATA[5], Q3_TXPLL_DRI_RDATA[4], 
        Q3_TXPLL_DRI_RDATA[3], Q3_TXPLL_DRI_RDATA[2], 
        Q3_TXPLL_DRI_RDATA[1], Q3_TXPLL_DRI_RDATA[0]}), 
        .Q3_TXPLL_DRI_INTERRUPT(Q3_TXPLL_DRI_INTERRUPT), 
        .Q5_TXPLL_DRI_CTRL({Q5_TXPLL_DRI_CTRL[10], 
        Q5_TXPLL_DRI_CTRL[9], Q5_TXPLL_DRI_CTRL[8], 
        Q5_TXPLL_DRI_CTRL[7], Q5_TXPLL_DRI_CTRL[6], 
        Q5_TXPLL_DRI_CTRL[5], Q5_TXPLL_DRI_CTRL[4], 
        Q5_TXPLL_DRI_CTRL[3], Q5_TXPLL_DRI_CTRL[2], 
        Q5_TXPLL_DRI_CTRL[1], Q5_TXPLL_DRI_CTRL[0]}), 
        .Q5_TXPLL_DRI_RDATA({Q5_TXPLL_DRI_RDATA[32], 
        Q5_TXPLL_DRI_RDATA[31], Q5_TXPLL_DRI_RDATA[30], 
        Q5_TXPLL_DRI_RDATA[29], Q5_TXPLL_DRI_RDATA[28], 
        Q5_TXPLL_DRI_RDATA[27], Q5_TXPLL_DRI_RDATA[26], 
        Q5_TXPLL_DRI_RDATA[25], Q5_TXPLL_DRI_RDATA[24], 
        Q5_TXPLL_DRI_RDATA[23], Q5_TXPLL_DRI_RDATA[22], 
        Q5_TXPLL_DRI_RDATA[21], Q5_TXPLL_DRI_RDATA[20], 
        Q5_TXPLL_DRI_RDATA[19], Q5_TXPLL_DRI_RDATA[18], 
        Q5_TXPLL_DRI_RDATA[17], Q5_TXPLL_DRI_RDATA[16], 
        Q5_TXPLL_DRI_RDATA[15], Q5_TXPLL_DRI_RDATA[14], 
        Q5_TXPLL_DRI_RDATA[13], Q5_TXPLL_DRI_RDATA[12], 
        Q5_TXPLL_DRI_RDATA[11], Q5_TXPLL_DRI_RDATA[10], 
        Q5_TXPLL_DRI_RDATA[9], Q5_TXPLL_DRI_RDATA[8], 
        Q5_TXPLL_DRI_RDATA[7], Q5_TXPLL_DRI_RDATA[6], 
        Q5_TXPLL_DRI_RDATA[5], Q5_TXPLL_DRI_RDATA[4], 
        Q5_TXPLL_DRI_RDATA[3], Q5_TXPLL_DRI_RDATA[2], 
        Q5_TXPLL_DRI_RDATA[1], Q5_TXPLL_DRI_RDATA[0]}), 
        .Q5_TXPLL_DRI_INTERRUPT(Q5_TXPLL_DRI_INTERRUPT), 
        .PLL0_NW_DRI_CTRL({PLL0_NW_DRI_CTRL[10], PLL0_NW_DRI_CTRL[9], 
        PLL0_NW_DRI_CTRL[8], PLL0_NW_DRI_CTRL[7], PLL0_NW_DRI_CTRL[6], 
        PLL0_NW_DRI_CTRL[5], PLL0_NW_DRI_CTRL[4], PLL0_NW_DRI_CTRL[3], 
        PLL0_NW_DRI_CTRL[2], PLL0_NW_DRI_CTRL[1], PLL0_NW_DRI_CTRL[0]})
        , .PLL0_NW_DRI_RDATA({PLL0_NW_DRI_RDATA[32], 
        PLL0_NW_DRI_RDATA[31], PLL0_NW_DRI_RDATA[30], 
        PLL0_NW_DRI_RDATA[29], PLL0_NW_DRI_RDATA[28], 
        PLL0_NW_DRI_RDATA[27], PLL0_NW_DRI_RDATA[26], 
        PLL0_NW_DRI_RDATA[25], PLL0_NW_DRI_RDATA[24], 
        PLL0_NW_DRI_RDATA[23], PLL0_NW_DRI_RDATA[22], 
        PLL0_NW_DRI_RDATA[21], PLL0_NW_DRI_RDATA[20], 
        PLL0_NW_DRI_RDATA[19], PLL0_NW_DRI_RDATA[18], 
        PLL0_NW_DRI_RDATA[17], PLL0_NW_DRI_RDATA[16], 
        PLL0_NW_DRI_RDATA[15], PLL0_NW_DRI_RDATA[14], 
        PLL0_NW_DRI_RDATA[13], PLL0_NW_DRI_RDATA[12], 
        PLL0_NW_DRI_RDATA[11], PLL0_NW_DRI_RDATA[10], 
        PLL0_NW_DRI_RDATA[9], PLL0_NW_DRI_RDATA[8], 
        PLL0_NW_DRI_RDATA[7], PLL0_NW_DRI_RDATA[6], 
        PLL0_NW_DRI_RDATA[5], PLL0_NW_DRI_RDATA[4], 
        PLL0_NW_DRI_RDATA[3], PLL0_NW_DRI_RDATA[2], 
        PLL0_NW_DRI_RDATA[1], PLL0_NW_DRI_RDATA[0]}), 
        .PLL0_NW_DRI_INTERRUPT(PLL0_NW_DRI_INTERRUPT), 
        .PLL1_NW_DRI_CTRL({PLL1_NW_DRI_CTRL[10], PLL1_NW_DRI_CTRL[9], 
        PLL1_NW_DRI_CTRL[8], PLL1_NW_DRI_CTRL[7], PLL1_NW_DRI_CTRL[6], 
        PLL1_NW_DRI_CTRL[5], PLL1_NW_DRI_CTRL[4], PLL1_NW_DRI_CTRL[3], 
        PLL1_NW_DRI_CTRL[2], PLL1_NW_DRI_CTRL[1], PLL1_NW_DRI_CTRL[0]})
        , .PLL1_NW_DRI_RDATA({PLL1_NW_DRI_RDATA[32], 
        PLL1_NW_DRI_RDATA[31], PLL1_NW_DRI_RDATA[30], 
        PLL1_NW_DRI_RDATA[29], PLL1_NW_DRI_RDATA[28], 
        PLL1_NW_DRI_RDATA[27], PLL1_NW_DRI_RDATA[26], 
        PLL1_NW_DRI_RDATA[25], PLL1_NW_DRI_RDATA[24], 
        PLL1_NW_DRI_RDATA[23], PLL1_NW_DRI_RDATA[22], 
        PLL1_NW_DRI_RDATA[21], PLL1_NW_DRI_RDATA[20], 
        PLL1_NW_DRI_RDATA[19], PLL1_NW_DRI_RDATA[18], 
        PLL1_NW_DRI_RDATA[17], PLL1_NW_DRI_RDATA[16], 
        PLL1_NW_DRI_RDATA[15], PLL1_NW_DRI_RDATA[14], 
        PLL1_NW_DRI_RDATA[13], PLL1_NW_DRI_RDATA[12], 
        PLL1_NW_DRI_RDATA[11], PLL1_NW_DRI_RDATA[10], 
        PLL1_NW_DRI_RDATA[9], PLL1_NW_DRI_RDATA[8], 
        PLL1_NW_DRI_RDATA[7], PLL1_NW_DRI_RDATA[6], 
        PLL1_NW_DRI_RDATA[5], PLL1_NW_DRI_RDATA[4], 
        PLL1_NW_DRI_RDATA[3], PLL1_NW_DRI_RDATA[2], 
        PLL1_NW_DRI_RDATA[1], PLL1_NW_DRI_RDATA[0]}), 
        .PLL1_NW_DRI_INTERRUPT(PLL1_NW_DRI_INTERRUPT), 
        .DLL0_NW_DRI_CTRL({DLL0_NW_DRI_CTRL[10], DLL0_NW_DRI_CTRL[9], 
        DLL0_NW_DRI_CTRL[8], DLL0_NW_DRI_CTRL[7], DLL0_NW_DRI_CTRL[6], 
        DLL0_NW_DRI_CTRL[5], DLL0_NW_DRI_CTRL[4], DLL0_NW_DRI_CTRL[3], 
        DLL0_NW_DRI_CTRL[2], DLL0_NW_DRI_CTRL[1], DLL0_NW_DRI_CTRL[0]})
        , .DLL0_NW_DRI_RDATA({DLL0_NW_DRI_RDATA[32], 
        DLL0_NW_DRI_RDATA[31], DLL0_NW_DRI_RDATA[30], 
        DLL0_NW_DRI_RDATA[29], DLL0_NW_DRI_RDATA[28], 
        DLL0_NW_DRI_RDATA[27], DLL0_NW_DRI_RDATA[26], 
        DLL0_NW_DRI_RDATA[25], DLL0_NW_DRI_RDATA[24], 
        DLL0_NW_DRI_RDATA[23], DLL0_NW_DRI_RDATA[22], 
        DLL0_NW_DRI_RDATA[21], DLL0_NW_DRI_RDATA[20], 
        DLL0_NW_DRI_RDATA[19], DLL0_NW_DRI_RDATA[18], 
        DLL0_NW_DRI_RDATA[17], DLL0_NW_DRI_RDATA[16], 
        DLL0_NW_DRI_RDATA[15], DLL0_NW_DRI_RDATA[14], 
        DLL0_NW_DRI_RDATA[13], DLL0_NW_DRI_RDATA[12], 
        DLL0_NW_DRI_RDATA[11], DLL0_NW_DRI_RDATA[10], 
        DLL0_NW_DRI_RDATA[9], DLL0_NW_DRI_RDATA[8], 
        DLL0_NW_DRI_RDATA[7], DLL0_NW_DRI_RDATA[6], 
        DLL0_NW_DRI_RDATA[5], DLL0_NW_DRI_RDATA[4], 
        DLL0_NW_DRI_RDATA[3], DLL0_NW_DRI_RDATA[2], 
        DLL0_NW_DRI_RDATA[1], DLL0_NW_DRI_RDATA[0]}), 
        .DLL0_NW_DRI_INTERRUPT(DLL0_NW_DRI_INTERRUPT), 
        .DLL1_NW_DRI_CTRL({DLL1_NW_DRI_CTRL[10], DLL1_NW_DRI_CTRL[9], 
        DLL1_NW_DRI_CTRL[8], DLL1_NW_DRI_CTRL[7], DLL1_NW_DRI_CTRL[6], 
        DLL1_NW_DRI_CTRL[5], DLL1_NW_DRI_CTRL[4], DLL1_NW_DRI_CTRL[3], 
        DLL1_NW_DRI_CTRL[2], DLL1_NW_DRI_CTRL[1], DLL1_NW_DRI_CTRL[0]})
        , .DLL1_NW_DRI_RDATA({DLL1_NW_DRI_RDATA[32], 
        DLL1_NW_DRI_RDATA[31], DLL1_NW_DRI_RDATA[30], 
        DLL1_NW_DRI_RDATA[29], DLL1_NW_DRI_RDATA[28], 
        DLL1_NW_DRI_RDATA[27], DLL1_NW_DRI_RDATA[26], 
        DLL1_NW_DRI_RDATA[25], DLL1_NW_DRI_RDATA[24], 
        DLL1_NW_DRI_RDATA[23], DLL1_NW_DRI_RDATA[22], 
        DLL1_NW_DRI_RDATA[21], DLL1_NW_DRI_RDATA[20], 
        DLL1_NW_DRI_RDATA[19], DLL1_NW_DRI_RDATA[18], 
        DLL1_NW_DRI_RDATA[17], DLL1_NW_DRI_RDATA[16], 
        DLL1_NW_DRI_RDATA[15], DLL1_NW_DRI_RDATA[14], 
        DLL1_NW_DRI_RDATA[13], DLL1_NW_DRI_RDATA[12], 
        DLL1_NW_DRI_RDATA[11], DLL1_NW_DRI_RDATA[10], 
        DLL1_NW_DRI_RDATA[9], DLL1_NW_DRI_RDATA[8], 
        DLL1_NW_DRI_RDATA[7], DLL1_NW_DRI_RDATA[6], 
        DLL1_NW_DRI_RDATA[5], DLL1_NW_DRI_RDATA[4], 
        DLL1_NW_DRI_RDATA[3], DLL1_NW_DRI_RDATA[2], 
        DLL1_NW_DRI_RDATA[1], DLL1_NW_DRI_RDATA[0]}), 
        .DLL1_NW_DRI_INTERRUPT(DLL1_NW_DRI_INTERRUPT), 
        .PLL0_NE_DRI_CTRL({PLL0_NE_DRI_CTRL[10], PLL0_NE_DRI_CTRL[9], 
        PLL0_NE_DRI_CTRL[8], PLL0_NE_DRI_CTRL[7], PLL0_NE_DRI_CTRL[6], 
        PLL0_NE_DRI_CTRL[5], PLL0_NE_DRI_CTRL[4], PLL0_NE_DRI_CTRL[3], 
        PLL0_NE_DRI_CTRL[2], PLL0_NE_DRI_CTRL[1], PLL0_NE_DRI_CTRL[0]})
        , .PLL0_NE_DRI_RDATA({PLL0_NE_DRI_RDATA[32], 
        PLL0_NE_DRI_RDATA[31], PLL0_NE_DRI_RDATA[30], 
        PLL0_NE_DRI_RDATA[29], PLL0_NE_DRI_RDATA[28], 
        PLL0_NE_DRI_RDATA[27], PLL0_NE_DRI_RDATA[26], 
        PLL0_NE_DRI_RDATA[25], PLL0_NE_DRI_RDATA[24], 
        PLL0_NE_DRI_RDATA[23], PLL0_NE_DRI_RDATA[22], 
        PLL0_NE_DRI_RDATA[21], PLL0_NE_DRI_RDATA[20], 
        PLL0_NE_DRI_RDATA[19], PLL0_NE_DRI_RDATA[18], 
        PLL0_NE_DRI_RDATA[17], PLL0_NE_DRI_RDATA[16], 
        PLL0_NE_DRI_RDATA[15], PLL0_NE_DRI_RDATA[14], 
        PLL0_NE_DRI_RDATA[13], PLL0_NE_DRI_RDATA[12], 
        PLL0_NE_DRI_RDATA[11], PLL0_NE_DRI_RDATA[10], 
        PLL0_NE_DRI_RDATA[9], PLL0_NE_DRI_RDATA[8], 
        PLL0_NE_DRI_RDATA[7], PLL0_NE_DRI_RDATA[6], 
        PLL0_NE_DRI_RDATA[5], PLL0_NE_DRI_RDATA[4], 
        PLL0_NE_DRI_RDATA[3], PLL0_NE_DRI_RDATA[2], 
        PLL0_NE_DRI_RDATA[1], PLL0_NE_DRI_RDATA[0]}), 
        .PLL0_NE_DRI_INTERRUPT(PLL0_NE_DRI_INTERRUPT), 
        .PLL1_NE_DRI_CTRL({PLL1_NE_DRI_CTRL[10], PLL1_NE_DRI_CTRL[9], 
        PLL1_NE_DRI_CTRL[8], PLL1_NE_DRI_CTRL[7], PLL1_NE_DRI_CTRL[6], 
        PLL1_NE_DRI_CTRL[5], PLL1_NE_DRI_CTRL[4], PLL1_NE_DRI_CTRL[3], 
        PLL1_NE_DRI_CTRL[2], PLL1_NE_DRI_CTRL[1], PLL1_NE_DRI_CTRL[0]})
        , .PLL1_NE_DRI_RDATA({PLL1_NE_DRI_RDATA[32], 
        PLL1_NE_DRI_RDATA[31], PLL1_NE_DRI_RDATA[30], 
        PLL1_NE_DRI_RDATA[29], PLL1_NE_DRI_RDATA[28], 
        PLL1_NE_DRI_RDATA[27], PLL1_NE_DRI_RDATA[26], 
        PLL1_NE_DRI_RDATA[25], PLL1_NE_DRI_RDATA[24], 
        PLL1_NE_DRI_RDATA[23], PLL1_NE_DRI_RDATA[22], 
        PLL1_NE_DRI_RDATA[21], PLL1_NE_DRI_RDATA[20], 
        PLL1_NE_DRI_RDATA[19], PLL1_NE_DRI_RDATA[18], 
        PLL1_NE_DRI_RDATA[17], PLL1_NE_DRI_RDATA[16], 
        PLL1_NE_DRI_RDATA[15], PLL1_NE_DRI_RDATA[14], 
        PLL1_NE_DRI_RDATA[13], PLL1_NE_DRI_RDATA[12], 
        PLL1_NE_DRI_RDATA[11], PLL1_NE_DRI_RDATA[10], 
        PLL1_NE_DRI_RDATA[9], PLL1_NE_DRI_RDATA[8], 
        PLL1_NE_DRI_RDATA[7], PLL1_NE_DRI_RDATA[6], 
        PLL1_NE_DRI_RDATA[5], PLL1_NE_DRI_RDATA[4], 
        PLL1_NE_DRI_RDATA[3], PLL1_NE_DRI_RDATA[2], 
        PLL1_NE_DRI_RDATA[1], PLL1_NE_DRI_RDATA[0]}), 
        .PLL1_NE_DRI_INTERRUPT(PLL1_NE_DRI_INTERRUPT), 
        .DLL0_NE_DRI_CTRL({DLL0_NE_DRI_CTRL[10], DLL0_NE_DRI_CTRL[9], 
        DLL0_NE_DRI_CTRL[8], DLL0_NE_DRI_CTRL[7], DLL0_NE_DRI_CTRL[6], 
        DLL0_NE_DRI_CTRL[5], DLL0_NE_DRI_CTRL[4], DLL0_NE_DRI_CTRL[3], 
        DLL0_NE_DRI_CTRL[2], DLL0_NE_DRI_CTRL[1], DLL0_NE_DRI_CTRL[0]})
        , .DLL0_NE_DRI_RDATA({DLL0_NE_DRI_RDATA[32], 
        DLL0_NE_DRI_RDATA[31], DLL0_NE_DRI_RDATA[30], 
        DLL0_NE_DRI_RDATA[29], DLL0_NE_DRI_RDATA[28], 
        DLL0_NE_DRI_RDATA[27], DLL0_NE_DRI_RDATA[26], 
        DLL0_NE_DRI_RDATA[25], DLL0_NE_DRI_RDATA[24], 
        DLL0_NE_DRI_RDATA[23], DLL0_NE_DRI_RDATA[22], 
        DLL0_NE_DRI_RDATA[21], DLL0_NE_DRI_RDATA[20], 
        DLL0_NE_DRI_RDATA[19], DLL0_NE_DRI_RDATA[18], 
        DLL0_NE_DRI_RDATA[17], DLL0_NE_DRI_RDATA[16], 
        DLL0_NE_DRI_RDATA[15], DLL0_NE_DRI_RDATA[14], 
        DLL0_NE_DRI_RDATA[13], DLL0_NE_DRI_RDATA[12], 
        DLL0_NE_DRI_RDATA[11], DLL0_NE_DRI_RDATA[10], 
        DLL0_NE_DRI_RDATA[9], DLL0_NE_DRI_RDATA[8], 
        DLL0_NE_DRI_RDATA[7], DLL0_NE_DRI_RDATA[6], 
        DLL0_NE_DRI_RDATA[5], DLL0_NE_DRI_RDATA[4], 
        DLL0_NE_DRI_RDATA[3], DLL0_NE_DRI_RDATA[2], 
        DLL0_NE_DRI_RDATA[1], DLL0_NE_DRI_RDATA[0]}), 
        .DLL0_NE_DRI_INTERRUPT(DLL0_NE_DRI_INTERRUPT), 
        .DLL1_NE_DRI_CTRL({DLL1_NE_DRI_CTRL[10], DLL1_NE_DRI_CTRL[9], 
        DLL1_NE_DRI_CTRL[8], DLL1_NE_DRI_CTRL[7], DLL1_NE_DRI_CTRL[6], 
        DLL1_NE_DRI_CTRL[5], DLL1_NE_DRI_CTRL[4], DLL1_NE_DRI_CTRL[3], 
        DLL1_NE_DRI_CTRL[2], DLL1_NE_DRI_CTRL[1], DLL1_NE_DRI_CTRL[0]})
        , .DLL1_NE_DRI_RDATA({DLL1_NE_DRI_RDATA[32], 
        DLL1_NE_DRI_RDATA[31], DLL1_NE_DRI_RDATA[30], 
        DLL1_NE_DRI_RDATA[29], DLL1_NE_DRI_RDATA[28], 
        DLL1_NE_DRI_RDATA[27], DLL1_NE_DRI_RDATA[26], 
        DLL1_NE_DRI_RDATA[25], DLL1_NE_DRI_RDATA[24], 
        DLL1_NE_DRI_RDATA[23], DLL1_NE_DRI_RDATA[22], 
        DLL1_NE_DRI_RDATA[21], DLL1_NE_DRI_RDATA[20], 
        DLL1_NE_DRI_RDATA[19], DLL1_NE_DRI_RDATA[18], 
        DLL1_NE_DRI_RDATA[17], DLL1_NE_DRI_RDATA[16], 
        DLL1_NE_DRI_RDATA[15], DLL1_NE_DRI_RDATA[14], 
        DLL1_NE_DRI_RDATA[13], DLL1_NE_DRI_RDATA[12], 
        DLL1_NE_DRI_RDATA[11], DLL1_NE_DRI_RDATA[10], 
        DLL1_NE_DRI_RDATA[9], DLL1_NE_DRI_RDATA[8], 
        DLL1_NE_DRI_RDATA[7], DLL1_NE_DRI_RDATA[6], 
        DLL1_NE_DRI_RDATA[5], DLL1_NE_DRI_RDATA[4], 
        DLL1_NE_DRI_RDATA[3], DLL1_NE_DRI_RDATA[2], 
        DLL1_NE_DRI_RDATA[1], DLL1_NE_DRI_RDATA[0]}), 
        .DLL1_NE_DRI_INTERRUPT(DLL1_NE_DRI_INTERRUPT), 
        .PLL0_SE_DRI_CTRL({PLL0_SE_DRI_CTRL[10], PLL0_SE_DRI_CTRL[9], 
        PLL0_SE_DRI_CTRL[8], PLL0_SE_DRI_CTRL[7], PLL0_SE_DRI_CTRL[6], 
        PLL0_SE_DRI_CTRL[5], PLL0_SE_DRI_CTRL[4], PLL0_SE_DRI_CTRL[3], 
        PLL0_SE_DRI_CTRL[2], PLL0_SE_DRI_CTRL[1], PLL0_SE_DRI_CTRL[0]})
        , .PLL0_SE_DRI_RDATA({PLL0_SE_DRI_RDATA[32], 
        PLL0_SE_DRI_RDATA[31], PLL0_SE_DRI_RDATA[30], 
        PLL0_SE_DRI_RDATA[29], PLL0_SE_DRI_RDATA[28], 
        PLL0_SE_DRI_RDATA[27], PLL0_SE_DRI_RDATA[26], 
        PLL0_SE_DRI_RDATA[25], PLL0_SE_DRI_RDATA[24], 
        PLL0_SE_DRI_RDATA[23], PLL0_SE_DRI_RDATA[22], 
        PLL0_SE_DRI_RDATA[21], PLL0_SE_DRI_RDATA[20], 
        PLL0_SE_DRI_RDATA[19], PLL0_SE_DRI_RDATA[18], 
        PLL0_SE_DRI_RDATA[17], PLL0_SE_DRI_RDATA[16], 
        PLL0_SE_DRI_RDATA[15], PLL0_SE_DRI_RDATA[14], 
        PLL0_SE_DRI_RDATA[13], PLL0_SE_DRI_RDATA[12], 
        PLL0_SE_DRI_RDATA[11], PLL0_SE_DRI_RDATA[10], 
        PLL0_SE_DRI_RDATA[9], PLL0_SE_DRI_RDATA[8], 
        PLL0_SE_DRI_RDATA[7], PLL0_SE_DRI_RDATA[6], 
        PLL0_SE_DRI_RDATA[5], PLL0_SE_DRI_RDATA[4], 
        PLL0_SE_DRI_RDATA[3], PLL0_SE_DRI_RDATA[2], 
        PLL0_SE_DRI_RDATA[1], PLL0_SE_DRI_RDATA[0]}), 
        .PLL0_SE_DRI_INTERRUPT(PLL0_SE_DRI_INTERRUPT), 
        .PLL1_SE_DRI_CTRL({PLL1_SE_DRI_CTRL[10], PLL1_SE_DRI_CTRL[9], 
        PLL1_SE_DRI_CTRL[8], PLL1_SE_DRI_CTRL[7], PLL1_SE_DRI_CTRL[6], 
        PLL1_SE_DRI_CTRL[5], PLL1_SE_DRI_CTRL[4], PLL1_SE_DRI_CTRL[3], 
        PLL1_SE_DRI_CTRL[2], PLL1_SE_DRI_CTRL[1], PLL1_SE_DRI_CTRL[0]})
        , .PLL1_SE_DRI_RDATA({PLL1_SE_DRI_RDATA[32], 
        PLL1_SE_DRI_RDATA[31], PLL1_SE_DRI_RDATA[30], 
        PLL1_SE_DRI_RDATA[29], PLL1_SE_DRI_RDATA[28], 
        PLL1_SE_DRI_RDATA[27], PLL1_SE_DRI_RDATA[26], 
        PLL1_SE_DRI_RDATA[25], PLL1_SE_DRI_RDATA[24], 
        PLL1_SE_DRI_RDATA[23], PLL1_SE_DRI_RDATA[22], 
        PLL1_SE_DRI_RDATA[21], PLL1_SE_DRI_RDATA[20], 
        PLL1_SE_DRI_RDATA[19], PLL1_SE_DRI_RDATA[18], 
        PLL1_SE_DRI_RDATA[17], PLL1_SE_DRI_RDATA[16], 
        PLL1_SE_DRI_RDATA[15], PLL1_SE_DRI_RDATA[14], 
        PLL1_SE_DRI_RDATA[13], PLL1_SE_DRI_RDATA[12], 
        PLL1_SE_DRI_RDATA[11], PLL1_SE_DRI_RDATA[10], 
        PLL1_SE_DRI_RDATA[9], PLL1_SE_DRI_RDATA[8], 
        PLL1_SE_DRI_RDATA[7], PLL1_SE_DRI_RDATA[6], 
        PLL1_SE_DRI_RDATA[5], PLL1_SE_DRI_RDATA[4], 
        PLL1_SE_DRI_RDATA[3], PLL1_SE_DRI_RDATA[2], 
        PLL1_SE_DRI_RDATA[1], PLL1_SE_DRI_RDATA[0]}), 
        .PLL1_SE_DRI_INTERRUPT(PLL1_SE_DRI_INTERRUPT), 
        .DLL0_SE_DRI_CTRL({DLL0_SE_DRI_CTRL[10], DLL0_SE_DRI_CTRL[9], 
        DLL0_SE_DRI_CTRL[8], DLL0_SE_DRI_CTRL[7], DLL0_SE_DRI_CTRL[6], 
        DLL0_SE_DRI_CTRL[5], DLL0_SE_DRI_CTRL[4], DLL0_SE_DRI_CTRL[3], 
        DLL0_SE_DRI_CTRL[2], DLL0_SE_DRI_CTRL[1], DLL0_SE_DRI_CTRL[0]})
        , .DLL0_SE_DRI_RDATA({DLL0_SE_DRI_RDATA[32], 
        DLL0_SE_DRI_RDATA[31], DLL0_SE_DRI_RDATA[30], 
        DLL0_SE_DRI_RDATA[29], DLL0_SE_DRI_RDATA[28], 
        DLL0_SE_DRI_RDATA[27], DLL0_SE_DRI_RDATA[26], 
        DLL0_SE_DRI_RDATA[25], DLL0_SE_DRI_RDATA[24], 
        DLL0_SE_DRI_RDATA[23], DLL0_SE_DRI_RDATA[22], 
        DLL0_SE_DRI_RDATA[21], DLL0_SE_DRI_RDATA[20], 
        DLL0_SE_DRI_RDATA[19], DLL0_SE_DRI_RDATA[18], 
        DLL0_SE_DRI_RDATA[17], DLL0_SE_DRI_RDATA[16], 
        DLL0_SE_DRI_RDATA[15], DLL0_SE_DRI_RDATA[14], 
        DLL0_SE_DRI_RDATA[13], DLL0_SE_DRI_RDATA[12], 
        DLL0_SE_DRI_RDATA[11], DLL0_SE_DRI_RDATA[10], 
        DLL0_SE_DRI_RDATA[9], DLL0_SE_DRI_RDATA[8], 
        DLL0_SE_DRI_RDATA[7], DLL0_SE_DRI_RDATA[6], 
        DLL0_SE_DRI_RDATA[5], DLL0_SE_DRI_RDATA[4], 
        DLL0_SE_DRI_RDATA[3], DLL0_SE_DRI_RDATA[2], 
        DLL0_SE_DRI_RDATA[1], DLL0_SE_DRI_RDATA[0]}), 
        .DLL0_SE_DRI_INTERRUPT(DLL0_SE_DRI_INTERRUPT), 
        .DLL1_SE_DRI_CTRL({DLL1_SE_DRI_CTRL[10], DLL1_SE_DRI_CTRL[9], 
        DLL1_SE_DRI_CTRL[8], DLL1_SE_DRI_CTRL[7], DLL1_SE_DRI_CTRL[6], 
        DLL1_SE_DRI_CTRL[5], DLL1_SE_DRI_CTRL[4], DLL1_SE_DRI_CTRL[3], 
        DLL1_SE_DRI_CTRL[2], DLL1_SE_DRI_CTRL[1], DLL1_SE_DRI_CTRL[0]})
        , .DLL1_SE_DRI_RDATA({DLL1_SE_DRI_RDATA[32], 
        DLL1_SE_DRI_RDATA[31], DLL1_SE_DRI_RDATA[30], 
        DLL1_SE_DRI_RDATA[29], DLL1_SE_DRI_RDATA[28], 
        DLL1_SE_DRI_RDATA[27], DLL1_SE_DRI_RDATA[26], 
        DLL1_SE_DRI_RDATA[25], DLL1_SE_DRI_RDATA[24], 
        DLL1_SE_DRI_RDATA[23], DLL1_SE_DRI_RDATA[22], 
        DLL1_SE_DRI_RDATA[21], DLL1_SE_DRI_RDATA[20], 
        DLL1_SE_DRI_RDATA[19], DLL1_SE_DRI_RDATA[18], 
        DLL1_SE_DRI_RDATA[17], DLL1_SE_DRI_RDATA[16], 
        DLL1_SE_DRI_RDATA[15], DLL1_SE_DRI_RDATA[14], 
        DLL1_SE_DRI_RDATA[13], DLL1_SE_DRI_RDATA[12], 
        DLL1_SE_DRI_RDATA[11], DLL1_SE_DRI_RDATA[10], 
        DLL1_SE_DRI_RDATA[9], DLL1_SE_DRI_RDATA[8], 
        DLL1_SE_DRI_RDATA[7], DLL1_SE_DRI_RDATA[6], 
        DLL1_SE_DRI_RDATA[5], DLL1_SE_DRI_RDATA[4], 
        DLL1_SE_DRI_RDATA[3], DLL1_SE_DRI_RDATA[2], 
        DLL1_SE_DRI_RDATA[1], DLL1_SE_DRI_RDATA[0]}), 
        .DLL1_SE_DRI_INTERRUPT(DLL1_SE_DRI_INTERRUPT), 
        .PLL0_SW_DRI_CTRL({PLL0_SW_DRI_CTRL[10], PLL0_SW_DRI_CTRL[9], 
        PLL0_SW_DRI_CTRL[8], PLL0_SW_DRI_CTRL[7], PLL0_SW_DRI_CTRL[6], 
        PLL0_SW_DRI_CTRL[5], PLL0_SW_DRI_CTRL[4], PLL0_SW_DRI_CTRL[3], 
        PLL0_SW_DRI_CTRL[2], PLL0_SW_DRI_CTRL[1], PLL0_SW_DRI_CTRL[0]})
        , .PLL0_SW_DRI_RDATA({PLL0_SW_DRI_RDATA[32], 
        PLL0_SW_DRI_RDATA[31], PLL0_SW_DRI_RDATA[30], 
        PLL0_SW_DRI_RDATA[29], PLL0_SW_DRI_RDATA[28], 
        PLL0_SW_DRI_RDATA[27], PLL0_SW_DRI_RDATA[26], 
        PLL0_SW_DRI_RDATA[25], PLL0_SW_DRI_RDATA[24], 
        PLL0_SW_DRI_RDATA[23], PLL0_SW_DRI_RDATA[22], 
        PLL0_SW_DRI_RDATA[21], PLL0_SW_DRI_RDATA[20], 
        PLL0_SW_DRI_RDATA[19], PLL0_SW_DRI_RDATA[18], 
        PLL0_SW_DRI_RDATA[17], PLL0_SW_DRI_RDATA[16], 
        PLL0_SW_DRI_RDATA[15], PLL0_SW_DRI_RDATA[14], 
        PLL0_SW_DRI_RDATA[13], PLL0_SW_DRI_RDATA[12], 
        PLL0_SW_DRI_RDATA[11], PLL0_SW_DRI_RDATA[10], 
        PLL0_SW_DRI_RDATA[9], PLL0_SW_DRI_RDATA[8], 
        PLL0_SW_DRI_RDATA[7], PLL0_SW_DRI_RDATA[6], 
        PLL0_SW_DRI_RDATA[5], PLL0_SW_DRI_RDATA[4], 
        PLL0_SW_DRI_RDATA[3], PLL0_SW_DRI_RDATA[2], 
        PLL0_SW_DRI_RDATA[1], PLL0_SW_DRI_RDATA[0]}), 
        .PLL0_SW_DRI_INTERRUPT(PLL0_SW_DRI_INTERRUPT), 
        .PLL1_SW_DRI_CTRL({PLL1_SW_DRI_CTRL[10], PLL1_SW_DRI_CTRL[9], 
        PLL1_SW_DRI_CTRL[8], PLL1_SW_DRI_CTRL[7], PLL1_SW_DRI_CTRL[6], 
        PLL1_SW_DRI_CTRL[5], PLL1_SW_DRI_CTRL[4], PLL1_SW_DRI_CTRL[3], 
        PLL1_SW_DRI_CTRL[2], PLL1_SW_DRI_CTRL[1], PLL1_SW_DRI_CTRL[0]})
        , .PLL1_SW_DRI_RDATA({PLL1_SW_DRI_RDATA[32], 
        PLL1_SW_DRI_RDATA[31], PLL1_SW_DRI_RDATA[30], 
        PLL1_SW_DRI_RDATA[29], PLL1_SW_DRI_RDATA[28], 
        PLL1_SW_DRI_RDATA[27], PLL1_SW_DRI_RDATA[26], 
        PLL1_SW_DRI_RDATA[25], PLL1_SW_DRI_RDATA[24], 
        PLL1_SW_DRI_RDATA[23], PLL1_SW_DRI_RDATA[22], 
        PLL1_SW_DRI_RDATA[21], PLL1_SW_DRI_RDATA[20], 
        PLL1_SW_DRI_RDATA[19], PLL1_SW_DRI_RDATA[18], 
        PLL1_SW_DRI_RDATA[17], PLL1_SW_DRI_RDATA[16], 
        PLL1_SW_DRI_RDATA[15], PLL1_SW_DRI_RDATA[14], 
        PLL1_SW_DRI_RDATA[13], PLL1_SW_DRI_RDATA[12], 
        PLL1_SW_DRI_RDATA[11], PLL1_SW_DRI_RDATA[10], 
        PLL1_SW_DRI_RDATA[9], PLL1_SW_DRI_RDATA[8], 
        PLL1_SW_DRI_RDATA[7], PLL1_SW_DRI_RDATA[6], 
        PLL1_SW_DRI_RDATA[5], PLL1_SW_DRI_RDATA[4], 
        PLL1_SW_DRI_RDATA[3], PLL1_SW_DRI_RDATA[2], 
        PLL1_SW_DRI_RDATA[1], PLL1_SW_DRI_RDATA[0]}), 
        .PLL1_SW_DRI_INTERRUPT(PLL1_SW_DRI_INTERRUPT), 
        .DLL0_SW_DRI_CTRL({DLL0_SW_DRI_CTRL[10], DLL0_SW_DRI_CTRL[9], 
        DLL0_SW_DRI_CTRL[8], DLL0_SW_DRI_CTRL[7], DLL0_SW_DRI_CTRL[6], 
        DLL0_SW_DRI_CTRL[5], DLL0_SW_DRI_CTRL[4], DLL0_SW_DRI_CTRL[3], 
        DLL0_SW_DRI_CTRL[2], DLL0_SW_DRI_CTRL[1], DLL0_SW_DRI_CTRL[0]})
        , .DLL0_SW_DRI_RDATA({DLL0_SW_DRI_RDATA[32], 
        DLL0_SW_DRI_RDATA[31], DLL0_SW_DRI_RDATA[30], 
        DLL0_SW_DRI_RDATA[29], DLL0_SW_DRI_RDATA[28], 
        DLL0_SW_DRI_RDATA[27], DLL0_SW_DRI_RDATA[26], 
        DLL0_SW_DRI_RDATA[25], DLL0_SW_DRI_RDATA[24], 
        DLL0_SW_DRI_RDATA[23], DLL0_SW_DRI_RDATA[22], 
        DLL0_SW_DRI_RDATA[21], DLL0_SW_DRI_RDATA[20], 
        DLL0_SW_DRI_RDATA[19], DLL0_SW_DRI_RDATA[18], 
        DLL0_SW_DRI_RDATA[17], DLL0_SW_DRI_RDATA[16], 
        DLL0_SW_DRI_RDATA[15], DLL0_SW_DRI_RDATA[14], 
        DLL0_SW_DRI_RDATA[13], DLL0_SW_DRI_RDATA[12], 
        DLL0_SW_DRI_RDATA[11], DLL0_SW_DRI_RDATA[10], 
        DLL0_SW_DRI_RDATA[9], DLL0_SW_DRI_RDATA[8], 
        DLL0_SW_DRI_RDATA[7], DLL0_SW_DRI_RDATA[6], 
        DLL0_SW_DRI_RDATA[5], DLL0_SW_DRI_RDATA[4], 
        DLL0_SW_DRI_RDATA[3], DLL0_SW_DRI_RDATA[2], 
        DLL0_SW_DRI_RDATA[1], DLL0_SW_DRI_RDATA[0]}), 
        .DLL0_SW_DRI_INTERRUPT(DLL0_SW_DRI_INTERRUPT), 
        .DLL1_SW_DRI_CTRL({DLL1_SW_DRI_CTRL[10], DLL1_SW_DRI_CTRL[9], 
        DLL1_SW_DRI_CTRL[8], DLL1_SW_DRI_CTRL[7], DLL1_SW_DRI_CTRL[6], 
        DLL1_SW_DRI_CTRL[5], DLL1_SW_DRI_CTRL[4], DLL1_SW_DRI_CTRL[3], 
        DLL1_SW_DRI_CTRL[2], DLL1_SW_DRI_CTRL[1], DLL1_SW_DRI_CTRL[0]})
        , .DLL1_SW_DRI_RDATA({DLL1_SW_DRI_RDATA[32], 
        DLL1_SW_DRI_RDATA[31], DLL1_SW_DRI_RDATA[30], 
        DLL1_SW_DRI_RDATA[29], DLL1_SW_DRI_RDATA[28], 
        DLL1_SW_DRI_RDATA[27], DLL1_SW_DRI_RDATA[26], 
        DLL1_SW_DRI_RDATA[25], DLL1_SW_DRI_RDATA[24], 
        DLL1_SW_DRI_RDATA[23], DLL1_SW_DRI_RDATA[22], 
        DLL1_SW_DRI_RDATA[21], DLL1_SW_DRI_RDATA[20], 
        DLL1_SW_DRI_RDATA[19], DLL1_SW_DRI_RDATA[18], 
        DLL1_SW_DRI_RDATA[17], DLL1_SW_DRI_RDATA[16], 
        DLL1_SW_DRI_RDATA[15], DLL1_SW_DRI_RDATA[14], 
        DLL1_SW_DRI_RDATA[13], DLL1_SW_DRI_RDATA[12], 
        DLL1_SW_DRI_RDATA[11], DLL1_SW_DRI_RDATA[10], 
        DLL1_SW_DRI_RDATA[9], DLL1_SW_DRI_RDATA[8], 
        DLL1_SW_DRI_RDATA[7], DLL1_SW_DRI_RDATA[6], 
        DLL1_SW_DRI_RDATA[5], DLL1_SW_DRI_RDATA[4], 
        DLL1_SW_DRI_RDATA[3], DLL1_SW_DRI_RDATA[2], 
        DLL1_SW_DRI_RDATA[1], DLL1_SW_DRI_RDATA[0]}), 
        .DLL1_SW_DRI_INTERRUPT(DLL1_SW_DRI_INTERRUPT), 
        .CRYPTO_DRI_CTRL({CRYPTO_DRI_CTRL[10], CRYPTO_DRI_CTRL[9], 
        CRYPTO_DRI_CTRL[8], CRYPTO_DRI_CTRL[7], CRYPTO_DRI_CTRL[6], 
        CRYPTO_DRI_CTRL[5], CRYPTO_DRI_CTRL[4], CRYPTO_DRI_CTRL[3], 
        CRYPTO_DRI_CTRL[2], CRYPTO_DRI_CTRL[1], CRYPTO_DRI_CTRL[0]}), 
        .CRYPTO_DRI_RDATA({CRYPTO_DRI_RDATA[32], CRYPTO_DRI_RDATA[31], 
        CRYPTO_DRI_RDATA[30], CRYPTO_DRI_RDATA[29], 
        CRYPTO_DRI_RDATA[28], CRYPTO_DRI_RDATA[27], 
        CRYPTO_DRI_RDATA[26], CRYPTO_DRI_RDATA[25], 
        CRYPTO_DRI_RDATA[24], CRYPTO_DRI_RDATA[23], 
        CRYPTO_DRI_RDATA[22], CRYPTO_DRI_RDATA[21], 
        CRYPTO_DRI_RDATA[20], CRYPTO_DRI_RDATA[19], 
        CRYPTO_DRI_RDATA[18], CRYPTO_DRI_RDATA[17], 
        CRYPTO_DRI_RDATA[16], CRYPTO_DRI_RDATA[15], 
        CRYPTO_DRI_RDATA[14], CRYPTO_DRI_RDATA[13], 
        CRYPTO_DRI_RDATA[12], CRYPTO_DRI_RDATA[11], 
        CRYPTO_DRI_RDATA[10], CRYPTO_DRI_RDATA[9], CRYPTO_DRI_RDATA[8], 
        CRYPTO_DRI_RDATA[7], CRYPTO_DRI_RDATA[6], CRYPTO_DRI_RDATA[5], 
        CRYPTO_DRI_RDATA[4], CRYPTO_DRI_RDATA[3], CRYPTO_DRI_RDATA[2], 
        CRYPTO_DRI_RDATA[1], CRYPTO_DRI_RDATA[0]}), 
        .CRYPTO_DRI_INTERRUPT(CRYPTO_DRI_INTERRUPT));
    
endmodule
